
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f8",x"ee",x"c2"),
    14 => (x"48",x"c4",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f1",x"e2"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"49",x"72"),
    82 => (x"c2",x"7c",x"71",x"99"),
    83 => (x"05",x"bf",x"c4",x"dc"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"c3",x"29",x"d8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"d0",x"49",x"66",x"d0"),
    90 => (x"99",x"ff",x"c3",x"29"),
    91 => (x"66",x"d0",x"7c",x"71"),
    92 => (x"c3",x"29",x"c8",x"49"),
    93 => (x"7c",x"71",x"99",x"ff"),
    94 => (x"c3",x"49",x"66",x"d0"),
    95 => (x"7c",x"71",x"99",x"ff"),
    96 => (x"29",x"d0",x"49",x"72"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"c9",x"4b",x"6c",x"7c"),
    99 => (x"c3",x"4d",x"ff",x"f0"),
   100 => (x"d0",x"05",x"ab",x"ff"),
   101 => (x"7c",x"ff",x"c3",x"87"),
   102 => (x"8d",x"c1",x"4b",x"6c"),
   103 => (x"c3",x"87",x"c6",x"02"),
   104 => (x"f0",x"02",x"ab",x"ff"),
   105 => (x"fe",x"48",x"73",x"87"),
   106 => (x"c0",x"1e",x"87",x"c7"),
   107 => (x"48",x"d4",x"ff",x"49"),
   108 => (x"c1",x"78",x"ff",x"c3"),
   109 => (x"b7",x"c8",x"c3",x"81"),
   110 => (x"87",x"f1",x"04",x"a9"),
   111 => (x"73",x"1e",x"4f",x"26"),
   112 => (x"c4",x"87",x"e7",x"1e"),
   113 => (x"c0",x"4b",x"df",x"f8"),
   114 => (x"f0",x"ff",x"c0",x"1e"),
   115 => (x"fd",x"49",x"f7",x"c1"),
   116 => (x"86",x"c4",x"87",x"e7"),
   117 => (x"c0",x"05",x"a8",x"c1"),
   118 => (x"d4",x"ff",x"87",x"ea"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"c0",x"c0",x"c0",x"c1"),
   121 => (x"c0",x"1e",x"c0",x"c0"),
   122 => (x"e9",x"c1",x"f0",x"e1"),
   123 => (x"87",x"c9",x"fd",x"49"),
   124 => (x"98",x"70",x"86",x"c4"),
   125 => (x"ff",x"87",x"ca",x"05"),
   126 => (x"ff",x"c3",x"48",x"d4"),
   127 => (x"cb",x"48",x"c1",x"78"),
   128 => (x"87",x"e6",x"fe",x"87"),
   129 => (x"fe",x"05",x"8b",x"c1"),
   130 => (x"48",x"c0",x"87",x"fd"),
   131 => (x"1e",x"87",x"e6",x"fc"),
   132 => (x"d4",x"ff",x"1e",x"73"),
   133 => (x"78",x"ff",x"c3",x"48"),
   134 => (x"1e",x"c0",x"4b",x"d3"),
   135 => (x"c1",x"f0",x"ff",x"c0"),
   136 => (x"d4",x"fc",x"49",x"c1"),
   137 => (x"70",x"86",x"c4",x"87"),
   138 => (x"87",x"ca",x"05",x"98"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"48",x"c1",x"78",x"ff"),
   141 => (x"f1",x"fd",x"87",x"cb"),
   142 => (x"05",x"8b",x"c1",x"87"),
   143 => (x"c0",x"87",x"db",x"ff"),
   144 => (x"87",x"f1",x"fb",x"48"),
   145 => (x"5c",x"5b",x"5e",x"0e"),
   146 => (x"4c",x"d4",x"ff",x"0e"),
   147 => (x"c6",x"87",x"db",x"fd"),
   148 => (x"e1",x"c0",x"1e",x"ea"),
   149 => (x"49",x"c8",x"c1",x"f0"),
   150 => (x"c4",x"87",x"de",x"fb"),
   151 => (x"02",x"a8",x"c1",x"86"),
   152 => (x"ea",x"fe",x"87",x"c8"),
   153 => (x"c1",x"48",x"c0",x"87"),
   154 => (x"da",x"fa",x"87",x"e2"),
   155 => (x"cf",x"49",x"70",x"87"),
   156 => (x"c6",x"99",x"ff",x"ff"),
   157 => (x"c8",x"02",x"a9",x"ea"),
   158 => (x"87",x"d3",x"fe",x"87"),
   159 => (x"cb",x"c1",x"48",x"c0"),
   160 => (x"7c",x"ff",x"c3",x"87"),
   161 => (x"fc",x"4b",x"f1",x"c0"),
   162 => (x"98",x"70",x"87",x"f4"),
   163 => (x"87",x"eb",x"c0",x"02"),
   164 => (x"ff",x"c0",x"1e",x"c0"),
   165 => (x"49",x"fa",x"c1",x"f0"),
   166 => (x"c4",x"87",x"de",x"fa"),
   167 => (x"05",x"98",x"70",x"86"),
   168 => (x"ff",x"c3",x"87",x"d9"),
   169 => (x"c3",x"49",x"6c",x"7c"),
   170 => (x"7c",x"7c",x"7c",x"ff"),
   171 => (x"99",x"c0",x"c1",x"7c"),
   172 => (x"c1",x"87",x"c4",x"02"),
   173 => (x"c0",x"87",x"d5",x"48"),
   174 => (x"c2",x"87",x"d1",x"48"),
   175 => (x"87",x"c4",x"05",x"ab"),
   176 => (x"87",x"c8",x"48",x"c0"),
   177 => (x"fe",x"05",x"8b",x"c1"),
   178 => (x"48",x"c0",x"87",x"fd"),
   179 => (x"1e",x"87",x"e4",x"f9"),
   180 => (x"dc",x"c2",x"1e",x"73"),
   181 => (x"78",x"c1",x"48",x"c4"),
   182 => (x"d0",x"ff",x"4b",x"c7"),
   183 => (x"fb",x"78",x"c2",x"48"),
   184 => (x"d0",x"ff",x"87",x"c8"),
   185 => (x"c0",x"78",x"c3",x"48"),
   186 => (x"d0",x"e5",x"c0",x"1e"),
   187 => (x"f9",x"49",x"c0",x"c1"),
   188 => (x"86",x"c4",x"87",x"c7"),
   189 => (x"c1",x"05",x"a8",x"c1"),
   190 => (x"ab",x"c2",x"4b",x"87"),
   191 => (x"c0",x"87",x"c5",x"05"),
   192 => (x"87",x"f9",x"c0",x"48"),
   193 => (x"ff",x"05",x"8b",x"c1"),
   194 => (x"f7",x"fc",x"87",x"d0"),
   195 => (x"c8",x"dc",x"c2",x"87"),
   196 => (x"05",x"98",x"70",x"58"),
   197 => (x"1e",x"c1",x"87",x"cd"),
   198 => (x"c1",x"f0",x"ff",x"c0"),
   199 => (x"d8",x"f8",x"49",x"d0"),
   200 => (x"ff",x"86",x"c4",x"87"),
   201 => (x"ff",x"c3",x"48",x"d4"),
   202 => (x"87",x"de",x"c4",x"78"),
   203 => (x"58",x"cc",x"dc",x"c2"),
   204 => (x"c2",x"48",x"d0",x"ff"),
   205 => (x"48",x"d4",x"ff",x"78"),
   206 => (x"c1",x"78",x"ff",x"c3"),
   207 => (x"87",x"f5",x"f7",x"48"),
   208 => (x"5c",x"5b",x"5e",x"0e"),
   209 => (x"4a",x"71",x"0e",x"5d"),
   210 => (x"ff",x"4d",x"ff",x"c3"),
   211 => (x"7c",x"75",x"4c",x"d4"),
   212 => (x"c4",x"48",x"d0",x"ff"),
   213 => (x"7c",x"75",x"78",x"c3"),
   214 => (x"ff",x"c0",x"1e",x"72"),
   215 => (x"49",x"d8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"d6",x"f7"),
   217 => (x"02",x"98",x"70",x"86"),
   218 => (x"48",x"c1",x"87",x"c5"),
   219 => (x"75",x"87",x"f0",x"c0"),
   220 => (x"7c",x"fe",x"c3",x"7c"),
   221 => (x"d4",x"1e",x"c0",x"c8"),
   222 => (x"fa",x"f4",x"49",x"66"),
   223 => (x"75",x"86",x"c4",x"87"),
   224 => (x"75",x"7c",x"75",x"7c"),
   225 => (x"e0",x"da",x"d8",x"7c"),
   226 => (x"6c",x"7c",x"75",x"4b"),
   227 => (x"c5",x"05",x"99",x"49"),
   228 => (x"05",x"8b",x"c1",x"87"),
   229 => (x"7c",x"75",x"87",x"f3"),
   230 => (x"c2",x"48",x"d0",x"ff"),
   231 => (x"f6",x"48",x"c0",x"78"),
   232 => (x"5e",x"0e",x"87",x"cf"),
   233 => (x"0e",x"5d",x"5c",x"5b"),
   234 => (x"4c",x"c0",x"4b",x"71"),
   235 => (x"df",x"cd",x"ee",x"c5"),
   236 => (x"48",x"d4",x"ff",x"4a"),
   237 => (x"68",x"78",x"ff",x"c3"),
   238 => (x"a9",x"fe",x"c3",x"49"),
   239 => (x"87",x"fd",x"c0",x"05"),
   240 => (x"9b",x"73",x"4d",x"70"),
   241 => (x"d0",x"87",x"cc",x"02"),
   242 => (x"49",x"73",x"1e",x"66"),
   243 => (x"c4",x"87",x"cf",x"f4"),
   244 => (x"ff",x"87",x"d6",x"86"),
   245 => (x"d1",x"c4",x"48",x"d0"),
   246 => (x"7d",x"ff",x"c3",x"78"),
   247 => (x"c1",x"48",x"66",x"d0"),
   248 => (x"58",x"a6",x"d4",x"88"),
   249 => (x"f0",x"05",x"98",x"70"),
   250 => (x"48",x"d4",x"ff",x"87"),
   251 => (x"78",x"78",x"ff",x"c3"),
   252 => (x"c5",x"05",x"9b",x"73"),
   253 => (x"48",x"d0",x"ff",x"87"),
   254 => (x"4a",x"c1",x"78",x"d0"),
   255 => (x"05",x"8a",x"c1",x"4c"),
   256 => (x"74",x"87",x"ee",x"fe"),
   257 => (x"87",x"e9",x"f4",x"48"),
   258 => (x"71",x"1e",x"73",x"1e"),
   259 => (x"ff",x"4b",x"c0",x"4a"),
   260 => (x"ff",x"c3",x"48",x"d4"),
   261 => (x"48",x"d0",x"ff",x"78"),
   262 => (x"ff",x"78",x"c3",x"c4"),
   263 => (x"ff",x"c3",x"48",x"d4"),
   264 => (x"c0",x"1e",x"72",x"78"),
   265 => (x"d1",x"c1",x"f0",x"ff"),
   266 => (x"87",x"cd",x"f4",x"49"),
   267 => (x"98",x"70",x"86",x"c4"),
   268 => (x"c8",x"87",x"d2",x"05"),
   269 => (x"66",x"cc",x"1e",x"c0"),
   270 => (x"87",x"e6",x"fd",x"49"),
   271 => (x"4b",x"70",x"86",x"c4"),
   272 => (x"c2",x"48",x"d0",x"ff"),
   273 => (x"f3",x"48",x"73",x"78"),
   274 => (x"5e",x"0e",x"87",x"eb"),
   275 => (x"0e",x"5d",x"5c",x"5b"),
   276 => (x"ff",x"c0",x"1e",x"c0"),
   277 => (x"49",x"c9",x"c1",x"f0"),
   278 => (x"d2",x"87",x"de",x"f3"),
   279 => (x"cc",x"dc",x"c2",x"1e"),
   280 => (x"87",x"fe",x"fc",x"49"),
   281 => (x"4c",x"c0",x"86",x"c8"),
   282 => (x"b7",x"d2",x"84",x"c1"),
   283 => (x"87",x"f8",x"04",x"ac"),
   284 => (x"97",x"cc",x"dc",x"c2"),
   285 => (x"c0",x"c3",x"49",x"bf"),
   286 => (x"a9",x"c0",x"c1",x"99"),
   287 => (x"87",x"e7",x"c0",x"05"),
   288 => (x"97",x"d3",x"dc",x"c2"),
   289 => (x"31",x"d0",x"49",x"bf"),
   290 => (x"97",x"d4",x"dc",x"c2"),
   291 => (x"32",x"c8",x"4a",x"bf"),
   292 => (x"dc",x"c2",x"b1",x"72"),
   293 => (x"4a",x"bf",x"97",x"d5"),
   294 => (x"cf",x"4c",x"71",x"b1"),
   295 => (x"9c",x"ff",x"ff",x"ff"),
   296 => (x"34",x"ca",x"84",x"c1"),
   297 => (x"c2",x"87",x"e7",x"c1"),
   298 => (x"bf",x"97",x"d5",x"dc"),
   299 => (x"c6",x"31",x"c1",x"49"),
   300 => (x"d6",x"dc",x"c2",x"99"),
   301 => (x"c7",x"4a",x"bf",x"97"),
   302 => (x"b1",x"72",x"2a",x"b7"),
   303 => (x"97",x"d1",x"dc",x"c2"),
   304 => (x"cf",x"4d",x"4a",x"bf"),
   305 => (x"d2",x"dc",x"c2",x"9d"),
   306 => (x"c3",x"4a",x"bf",x"97"),
   307 => (x"c2",x"32",x"ca",x"9a"),
   308 => (x"bf",x"97",x"d3",x"dc"),
   309 => (x"73",x"33",x"c2",x"4b"),
   310 => (x"d4",x"dc",x"c2",x"b2"),
   311 => (x"c3",x"4b",x"bf",x"97"),
   312 => (x"b7",x"c6",x"9b",x"c0"),
   313 => (x"c2",x"b2",x"73",x"2b"),
   314 => (x"71",x"48",x"c1",x"81"),
   315 => (x"c1",x"49",x"70",x"30"),
   316 => (x"70",x"30",x"75",x"48"),
   317 => (x"c1",x"4c",x"72",x"4d"),
   318 => (x"c8",x"94",x"71",x"84"),
   319 => (x"06",x"ad",x"b7",x"c0"),
   320 => (x"34",x"c1",x"87",x"cc"),
   321 => (x"c0",x"c8",x"2d",x"b7"),
   322 => (x"ff",x"01",x"ad",x"b7"),
   323 => (x"48",x"74",x"87",x"f4"),
   324 => (x"0e",x"87",x"de",x"f0"),
   325 => (x"5d",x"5c",x"5b",x"5e"),
   326 => (x"c2",x"86",x"f8",x"0e"),
   327 => (x"c0",x"48",x"f2",x"e4"),
   328 => (x"ea",x"dc",x"c2",x"78"),
   329 => (x"fb",x"49",x"c0",x"1e"),
   330 => (x"86",x"c4",x"87",x"de"),
   331 => (x"c5",x"05",x"98",x"70"),
   332 => (x"c9",x"48",x"c0",x"87"),
   333 => (x"4d",x"c0",x"87",x"ce"),
   334 => (x"f2",x"c0",x"7e",x"c1"),
   335 => (x"c2",x"49",x"bf",x"ec"),
   336 => (x"71",x"4a",x"e0",x"dd"),
   337 => (x"e0",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"7e",x"c0",x"87",x"c2"),
   340 => (x"bf",x"e8",x"f2",x"c0"),
   341 => (x"fc",x"dd",x"c2",x"49"),
   342 => (x"4b",x"c8",x"71",x"4a"),
   343 => (x"70",x"87",x"ca",x"ec"),
   344 => (x"87",x"c2",x"05",x"98"),
   345 => (x"02",x"6e",x"7e",x"c0"),
   346 => (x"c2",x"87",x"fd",x"c0"),
   347 => (x"4d",x"bf",x"f0",x"e3"),
   348 => (x"9f",x"e8",x"e4",x"c2"),
   349 => (x"c5",x"48",x"7e",x"bf"),
   350 => (x"05",x"a8",x"ea",x"d6"),
   351 => (x"e3",x"c2",x"87",x"c7"),
   352 => (x"ce",x"4d",x"bf",x"f0"),
   353 => (x"ca",x"48",x"6e",x"87"),
   354 => (x"02",x"a8",x"d5",x"e9"),
   355 => (x"48",x"c0",x"87",x"c5"),
   356 => (x"c2",x"87",x"f1",x"c7"),
   357 => (x"75",x"1e",x"ea",x"dc"),
   358 => (x"87",x"ec",x"f9",x"49"),
   359 => (x"98",x"70",x"86",x"c4"),
   360 => (x"c0",x"87",x"c5",x"05"),
   361 => (x"87",x"dc",x"c7",x"48"),
   362 => (x"bf",x"e8",x"f2",x"c0"),
   363 => (x"fc",x"dd",x"c2",x"49"),
   364 => (x"4b",x"c8",x"71",x"4a"),
   365 => (x"70",x"87",x"f2",x"ea"),
   366 => (x"87",x"c8",x"05",x"98"),
   367 => (x"48",x"f2",x"e4",x"c2"),
   368 => (x"87",x"da",x"78",x"c1"),
   369 => (x"bf",x"ec",x"f2",x"c0"),
   370 => (x"e0",x"dd",x"c2",x"49"),
   371 => (x"4b",x"c8",x"71",x"4a"),
   372 => (x"70",x"87",x"d6",x"ea"),
   373 => (x"c5",x"c0",x"02",x"98"),
   374 => (x"c6",x"48",x"c0",x"87"),
   375 => (x"e4",x"c2",x"87",x"e6"),
   376 => (x"49",x"bf",x"97",x"e8"),
   377 => (x"05",x"a9",x"d5",x"c1"),
   378 => (x"c2",x"87",x"cd",x"c0"),
   379 => (x"bf",x"97",x"e9",x"e4"),
   380 => (x"a9",x"ea",x"c2",x"49"),
   381 => (x"87",x"c5",x"c0",x"02"),
   382 => (x"c7",x"c6",x"48",x"c0"),
   383 => (x"ea",x"dc",x"c2",x"87"),
   384 => (x"48",x"7e",x"bf",x"97"),
   385 => (x"02",x"a8",x"e9",x"c3"),
   386 => (x"6e",x"87",x"ce",x"c0"),
   387 => (x"a8",x"eb",x"c3",x"48"),
   388 => (x"87",x"c5",x"c0",x"02"),
   389 => (x"eb",x"c5",x"48",x"c0"),
   390 => (x"f5",x"dc",x"c2",x"87"),
   391 => (x"99",x"49",x"bf",x"97"),
   392 => (x"87",x"cc",x"c0",x"05"),
   393 => (x"97",x"f6",x"dc",x"c2"),
   394 => (x"a9",x"c2",x"49",x"bf"),
   395 => (x"87",x"c5",x"c0",x"02"),
   396 => (x"cf",x"c5",x"48",x"c0"),
   397 => (x"f7",x"dc",x"c2",x"87"),
   398 => (x"c2",x"48",x"bf",x"97"),
   399 => (x"70",x"58",x"ee",x"e4"),
   400 => (x"88",x"c1",x"48",x"4c"),
   401 => (x"58",x"f2",x"e4",x"c2"),
   402 => (x"97",x"f8",x"dc",x"c2"),
   403 => (x"81",x"75",x"49",x"bf"),
   404 => (x"97",x"f9",x"dc",x"c2"),
   405 => (x"32",x"c8",x"4a",x"bf"),
   406 => (x"c2",x"7e",x"a1",x"72"),
   407 => (x"6e",x"48",x"ff",x"e8"),
   408 => (x"fa",x"dc",x"c2",x"78"),
   409 => (x"c8",x"48",x"bf",x"97"),
   410 => (x"e4",x"c2",x"58",x"a6"),
   411 => (x"c2",x"02",x"bf",x"f2"),
   412 => (x"f2",x"c0",x"87",x"d4"),
   413 => (x"c2",x"49",x"bf",x"e8"),
   414 => (x"71",x"4a",x"fc",x"dd"),
   415 => (x"e8",x"e7",x"4b",x"c8"),
   416 => (x"02",x"98",x"70",x"87"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"f8",x"c3",x"48"),
   419 => (x"bf",x"ea",x"e4",x"c2"),
   420 => (x"d3",x"e9",x"c2",x"4c"),
   421 => (x"cf",x"dd",x"c2",x"5c"),
   422 => (x"c8",x"49",x"bf",x"97"),
   423 => (x"ce",x"dd",x"c2",x"31"),
   424 => (x"a1",x"4a",x"bf",x"97"),
   425 => (x"d0",x"dd",x"c2",x"49"),
   426 => (x"d0",x"4a",x"bf",x"97"),
   427 => (x"49",x"a1",x"72",x"32"),
   428 => (x"97",x"d1",x"dd",x"c2"),
   429 => (x"32",x"d8",x"4a",x"bf"),
   430 => (x"c4",x"49",x"a1",x"72"),
   431 => (x"e8",x"c2",x"91",x"66"),
   432 => (x"c2",x"81",x"bf",x"ff"),
   433 => (x"c2",x"59",x"c7",x"e9"),
   434 => (x"bf",x"97",x"d7",x"dd"),
   435 => (x"c2",x"32",x"c8",x"4a"),
   436 => (x"bf",x"97",x"d6",x"dd"),
   437 => (x"c2",x"4a",x"a2",x"4b"),
   438 => (x"bf",x"97",x"d8",x"dd"),
   439 => (x"73",x"33",x"d0",x"4b"),
   440 => (x"dd",x"c2",x"4a",x"a2"),
   441 => (x"4b",x"bf",x"97",x"d9"),
   442 => (x"33",x"d8",x"9b",x"cf"),
   443 => (x"c2",x"4a",x"a2",x"73"),
   444 => (x"c2",x"5a",x"cb",x"e9"),
   445 => (x"4a",x"bf",x"c7",x"e9"),
   446 => (x"92",x"74",x"8a",x"c2"),
   447 => (x"48",x"cb",x"e9",x"c2"),
   448 => (x"c1",x"78",x"a1",x"72"),
   449 => (x"dc",x"c2",x"87",x"ca"),
   450 => (x"49",x"bf",x"97",x"fc"),
   451 => (x"dc",x"c2",x"31",x"c8"),
   452 => (x"4a",x"bf",x"97",x"fb"),
   453 => (x"e4",x"c2",x"49",x"a1"),
   454 => (x"e4",x"c2",x"59",x"fa"),
   455 => (x"c5",x"49",x"bf",x"f6"),
   456 => (x"81",x"ff",x"c7",x"31"),
   457 => (x"e9",x"c2",x"29",x"c9"),
   458 => (x"dd",x"c2",x"59",x"d3"),
   459 => (x"4a",x"bf",x"97",x"c1"),
   460 => (x"dd",x"c2",x"32",x"c8"),
   461 => (x"4b",x"bf",x"97",x"c0"),
   462 => (x"66",x"c4",x"4a",x"a2"),
   463 => (x"c2",x"82",x"6e",x"92"),
   464 => (x"c2",x"5a",x"cf",x"e9"),
   465 => (x"c0",x"48",x"c7",x"e9"),
   466 => (x"c3",x"e9",x"c2",x"78"),
   467 => (x"78",x"a1",x"72",x"48"),
   468 => (x"48",x"d3",x"e9",x"c2"),
   469 => (x"bf",x"c7",x"e9",x"c2"),
   470 => (x"d7",x"e9",x"c2",x"78"),
   471 => (x"cb",x"e9",x"c2",x"48"),
   472 => (x"e4",x"c2",x"78",x"bf"),
   473 => (x"c0",x"02",x"bf",x"f2"),
   474 => (x"48",x"74",x"87",x"c9"),
   475 => (x"7e",x"70",x"30",x"c4"),
   476 => (x"c2",x"87",x"c9",x"c0"),
   477 => (x"48",x"bf",x"cf",x"e9"),
   478 => (x"7e",x"70",x"30",x"c4"),
   479 => (x"48",x"f6",x"e4",x"c2"),
   480 => (x"48",x"c1",x"78",x"6e"),
   481 => (x"4d",x"26",x"8e",x"f8"),
   482 => (x"4b",x"26",x"4c",x"26"),
   483 => (x"5e",x"0e",x"4f",x"26"),
   484 => (x"0e",x"5d",x"5c",x"5b"),
   485 => (x"e4",x"c2",x"4a",x"71"),
   486 => (x"cb",x"02",x"bf",x"f2"),
   487 => (x"c7",x"4b",x"72",x"87"),
   488 => (x"c1",x"4c",x"72",x"2b"),
   489 => (x"87",x"c9",x"9c",x"ff"),
   490 => (x"2b",x"c8",x"4b",x"72"),
   491 => (x"ff",x"c3",x"4c",x"72"),
   492 => (x"ff",x"e8",x"c2",x"9c"),
   493 => (x"f2",x"c0",x"83",x"bf"),
   494 => (x"02",x"ab",x"bf",x"e4"),
   495 => (x"f2",x"c0",x"87",x"d9"),
   496 => (x"dc",x"c2",x"5b",x"e8"),
   497 => (x"49",x"73",x"1e",x"ea"),
   498 => (x"c4",x"87",x"fd",x"f0"),
   499 => (x"05",x"98",x"70",x"86"),
   500 => (x"48",x"c0",x"87",x"c5"),
   501 => (x"c2",x"87",x"e6",x"c0"),
   502 => (x"02",x"bf",x"f2",x"e4"),
   503 => (x"49",x"74",x"87",x"d2"),
   504 => (x"dc",x"c2",x"91",x"c4"),
   505 => (x"4d",x"69",x"81",x"ea"),
   506 => (x"ff",x"ff",x"ff",x"cf"),
   507 => (x"87",x"cb",x"9d",x"ff"),
   508 => (x"91",x"c2",x"49",x"74"),
   509 => (x"81",x"ea",x"dc",x"c2"),
   510 => (x"75",x"4d",x"69",x"9f"),
   511 => (x"87",x"c6",x"fe",x"48"),
   512 => (x"5c",x"5b",x"5e",x"0e"),
   513 => (x"86",x"f8",x"0e",x"5d"),
   514 => (x"05",x"9c",x"4c",x"71"),
   515 => (x"48",x"c0",x"87",x"c5"),
   516 => (x"c8",x"87",x"c1",x"c3"),
   517 => (x"c0",x"48",x"7e",x"a4"),
   518 => (x"02",x"66",x"d8",x"78"),
   519 => (x"66",x"d8",x"87",x"c7"),
   520 => (x"c5",x"05",x"bf",x"97"),
   521 => (x"c2",x"48",x"c0",x"87"),
   522 => (x"1e",x"c0",x"87",x"ea"),
   523 => (x"ca",x"49",x"49",x"c1"),
   524 => (x"86",x"c4",x"87",x"d7"),
   525 => (x"02",x"9d",x"4d",x"70"),
   526 => (x"c2",x"87",x"c2",x"c1"),
   527 => (x"d8",x"4a",x"fa",x"e4"),
   528 => (x"c9",x"e0",x"49",x"66"),
   529 => (x"02",x"98",x"70",x"87"),
   530 => (x"75",x"87",x"f2",x"c0"),
   531 => (x"49",x"66",x"d8",x"4a"),
   532 => (x"ee",x"e0",x"4b",x"cb"),
   533 => (x"02",x"98",x"70",x"87"),
   534 => (x"c0",x"87",x"e2",x"c0"),
   535 => (x"02",x"9d",x"75",x"1e"),
   536 => (x"a6",x"c8",x"87",x"c7"),
   537 => (x"c5",x"78",x"c0",x"48"),
   538 => (x"48",x"a6",x"c8",x"87"),
   539 => (x"66",x"c8",x"78",x"c1"),
   540 => (x"87",x"d5",x"c9",x"49"),
   541 => (x"4d",x"70",x"86",x"c4"),
   542 => (x"fe",x"fe",x"05",x"9d"),
   543 => (x"02",x"9d",x"75",x"87"),
   544 => (x"dc",x"87",x"cf",x"c1"),
   545 => (x"48",x"6e",x"49",x"a5"),
   546 => (x"a5",x"da",x"78",x"69"),
   547 => (x"48",x"a6",x"c4",x"49"),
   548 => (x"9f",x"78",x"a4",x"c4"),
   549 => (x"66",x"c4",x"48",x"69"),
   550 => (x"e4",x"c2",x"78",x"08"),
   551 => (x"d2",x"02",x"bf",x"f2"),
   552 => (x"49",x"a5",x"d4",x"87"),
   553 => (x"c0",x"49",x"69",x"9f"),
   554 => (x"71",x"99",x"ff",x"ff"),
   555 => (x"70",x"30",x"d0",x"48"),
   556 => (x"c0",x"87",x"c2",x"7e"),
   557 => (x"48",x"49",x"6e",x"7e"),
   558 => (x"80",x"bf",x"66",x"c4"),
   559 => (x"78",x"08",x"66",x"c4"),
   560 => (x"a4",x"cc",x"7c",x"c0"),
   561 => (x"bf",x"66",x"c4",x"49"),
   562 => (x"49",x"a4",x"d0",x"79"),
   563 => (x"48",x"c1",x"79",x"c0"),
   564 => (x"48",x"c0",x"87",x"c2"),
   565 => (x"ed",x"fa",x"8e",x"f8"),
   566 => (x"5b",x"5e",x"0e",x"87"),
   567 => (x"71",x"0e",x"5d",x"5c"),
   568 => (x"c1",x"02",x"9c",x"4c"),
   569 => (x"a4",x"c8",x"87",x"ca"),
   570 => (x"c1",x"02",x"69",x"49"),
   571 => (x"66",x"d0",x"87",x"c2"),
   572 => (x"82",x"49",x"6c",x"4a"),
   573 => (x"d0",x"5a",x"a6",x"d4"),
   574 => (x"c2",x"b9",x"4d",x"66"),
   575 => (x"4a",x"bf",x"ee",x"e4"),
   576 => (x"99",x"72",x"ba",x"ff"),
   577 => (x"c0",x"02",x"99",x"71"),
   578 => (x"a4",x"c4",x"87",x"e4"),
   579 => (x"f9",x"49",x"6b",x"4b"),
   580 => (x"7b",x"70",x"87",x"fc"),
   581 => (x"bf",x"ea",x"e4",x"c2"),
   582 => (x"71",x"81",x"6c",x"49"),
   583 => (x"c2",x"b9",x"75",x"7c"),
   584 => (x"4a",x"bf",x"ee",x"e4"),
   585 => (x"99",x"72",x"ba",x"ff"),
   586 => (x"ff",x"05",x"99",x"71"),
   587 => (x"7c",x"75",x"87",x"dc"),
   588 => (x"1e",x"87",x"d3",x"f9"),
   589 => (x"4b",x"71",x"1e",x"73"),
   590 => (x"87",x"c7",x"02",x"9b"),
   591 => (x"69",x"49",x"a3",x"c8"),
   592 => (x"c0",x"87",x"c5",x"05"),
   593 => (x"87",x"f7",x"c0",x"48"),
   594 => (x"bf",x"c3",x"e9",x"c2"),
   595 => (x"49",x"a3",x"c4",x"4a"),
   596 => (x"89",x"c2",x"49",x"69"),
   597 => (x"bf",x"ea",x"e4",x"c2"),
   598 => (x"4a",x"a2",x"71",x"91"),
   599 => (x"bf",x"ee",x"e4",x"c2"),
   600 => (x"71",x"99",x"6b",x"49"),
   601 => (x"f2",x"c0",x"4a",x"a2"),
   602 => (x"66",x"c8",x"5a",x"e8"),
   603 => (x"ea",x"49",x"72",x"1e"),
   604 => (x"86",x"c4",x"87",x"d6"),
   605 => (x"c4",x"05",x"98",x"70"),
   606 => (x"c2",x"48",x"c0",x"87"),
   607 => (x"f8",x"48",x"c1",x"87"),
   608 => (x"73",x"1e",x"87",x"c8"),
   609 => (x"9b",x"4b",x"71",x"1e"),
   610 => (x"c8",x"87",x"c7",x"02"),
   611 => (x"05",x"69",x"49",x"a3"),
   612 => (x"48",x"c0",x"87",x"c5"),
   613 => (x"c2",x"87",x"f7",x"c0"),
   614 => (x"4a",x"bf",x"c3",x"e9"),
   615 => (x"69",x"49",x"a3",x"c4"),
   616 => (x"c2",x"89",x"c2",x"49"),
   617 => (x"91",x"bf",x"ea",x"e4"),
   618 => (x"c2",x"4a",x"a2",x"71"),
   619 => (x"49",x"bf",x"ee",x"e4"),
   620 => (x"a2",x"71",x"99",x"6b"),
   621 => (x"e8",x"f2",x"c0",x"4a"),
   622 => (x"1e",x"66",x"c8",x"5a"),
   623 => (x"ff",x"e5",x"49",x"72"),
   624 => (x"70",x"86",x"c4",x"87"),
   625 => (x"87",x"c4",x"05",x"98"),
   626 => (x"87",x"c2",x"48",x"c0"),
   627 => (x"f9",x"f6",x"48",x"c1"),
   628 => (x"5b",x"5e",x"0e",x"87"),
   629 => (x"1e",x"0e",x"5d",x"5c"),
   630 => (x"66",x"d4",x"4b",x"71"),
   631 => (x"02",x"9b",x"73",x"4d"),
   632 => (x"c8",x"87",x"cc",x"c1"),
   633 => (x"02",x"69",x"49",x"a3"),
   634 => (x"d0",x"87",x"c4",x"c1"),
   635 => (x"e4",x"c2",x"4c",x"a3"),
   636 => (x"ff",x"49",x"bf",x"ee"),
   637 => (x"99",x"4a",x"6c",x"b9"),
   638 => (x"a9",x"66",x"d4",x"7e"),
   639 => (x"c0",x"87",x"cd",x"06"),
   640 => (x"a3",x"cc",x"7c",x"7b"),
   641 => (x"49",x"a3",x"c4",x"4a"),
   642 => (x"87",x"ca",x"79",x"6a"),
   643 => (x"c0",x"f8",x"49",x"72"),
   644 => (x"4d",x"66",x"d4",x"99"),
   645 => (x"49",x"75",x"8d",x"71"),
   646 => (x"1e",x"71",x"29",x"c9"),
   647 => (x"f8",x"fa",x"49",x"73"),
   648 => (x"ea",x"dc",x"c2",x"87"),
   649 => (x"fc",x"49",x"73",x"1e"),
   650 => (x"86",x"c8",x"87",x"c9"),
   651 => (x"26",x"7c",x"66",x"d4"),
   652 => (x"1e",x"87",x"d3",x"f5"),
   653 => (x"4b",x"71",x"1e",x"73"),
   654 => (x"e4",x"c0",x"02",x"9b"),
   655 => (x"d7",x"e9",x"c2",x"87"),
   656 => (x"c2",x"4a",x"73",x"5b"),
   657 => (x"ea",x"e4",x"c2",x"8a"),
   658 => (x"c2",x"92",x"49",x"bf"),
   659 => (x"48",x"bf",x"c3",x"e9"),
   660 => (x"e9",x"c2",x"80",x"72"),
   661 => (x"48",x"71",x"58",x"db"),
   662 => (x"e4",x"c2",x"30",x"c4"),
   663 => (x"ed",x"c0",x"58",x"fa"),
   664 => (x"d3",x"e9",x"c2",x"87"),
   665 => (x"c7",x"e9",x"c2",x"48"),
   666 => (x"e9",x"c2",x"78",x"bf"),
   667 => (x"e9",x"c2",x"48",x"d7"),
   668 => (x"c2",x"78",x"bf",x"cb"),
   669 => (x"02",x"bf",x"f2",x"e4"),
   670 => (x"e4",x"c2",x"87",x"c9"),
   671 => (x"c4",x"49",x"bf",x"ea"),
   672 => (x"c2",x"87",x"c7",x"31"),
   673 => (x"49",x"bf",x"cf",x"e9"),
   674 => (x"e4",x"c2",x"31",x"c4"),
   675 => (x"f9",x"f3",x"59",x"fa"),
   676 => (x"5b",x"5e",x"0e",x"87"),
   677 => (x"4a",x"71",x"0e",x"5c"),
   678 => (x"9a",x"72",x"4b",x"c0"),
   679 => (x"87",x"e1",x"c0",x"02"),
   680 => (x"9f",x"49",x"a2",x"da"),
   681 => (x"e4",x"c2",x"4b",x"69"),
   682 => (x"cf",x"02",x"bf",x"f2"),
   683 => (x"49",x"a2",x"d4",x"87"),
   684 => (x"4c",x"49",x"69",x"9f"),
   685 => (x"9c",x"ff",x"ff",x"c0"),
   686 => (x"87",x"c2",x"34",x"d0"),
   687 => (x"49",x"74",x"4c",x"c0"),
   688 => (x"fd",x"49",x"73",x"b3"),
   689 => (x"ff",x"f2",x"87",x"ed"),
   690 => (x"5b",x"5e",x"0e",x"87"),
   691 => (x"f4",x"0e",x"5d",x"5c"),
   692 => (x"c0",x"4a",x"71",x"86"),
   693 => (x"02",x"9a",x"72",x"7e"),
   694 => (x"dc",x"c2",x"87",x"d8"),
   695 => (x"78",x"c0",x"48",x"e6"),
   696 => (x"48",x"de",x"dc",x"c2"),
   697 => (x"bf",x"d7",x"e9",x"c2"),
   698 => (x"e2",x"dc",x"c2",x"78"),
   699 => (x"d3",x"e9",x"c2",x"48"),
   700 => (x"e5",x"c2",x"78",x"bf"),
   701 => (x"50",x"c0",x"48",x"c7"),
   702 => (x"bf",x"f6",x"e4",x"c2"),
   703 => (x"e6",x"dc",x"c2",x"49"),
   704 => (x"aa",x"71",x"4a",x"bf"),
   705 => (x"87",x"c9",x"c4",x"03"),
   706 => (x"99",x"cf",x"49",x"72"),
   707 => (x"87",x"e9",x"c0",x"05"),
   708 => (x"48",x"e4",x"f2",x"c0"),
   709 => (x"bf",x"de",x"dc",x"c2"),
   710 => (x"ea",x"dc",x"c2",x"78"),
   711 => (x"de",x"dc",x"c2",x"1e"),
   712 => (x"dc",x"c2",x"49",x"bf"),
   713 => (x"a1",x"c1",x"48",x"de"),
   714 => (x"db",x"e3",x"71",x"78"),
   715 => (x"c0",x"86",x"c4",x"87"),
   716 => (x"c2",x"48",x"e0",x"f2"),
   717 => (x"cc",x"78",x"ea",x"dc"),
   718 => (x"e0",x"f2",x"c0",x"87"),
   719 => (x"e0",x"c0",x"48",x"bf"),
   720 => (x"e4",x"f2",x"c0",x"80"),
   721 => (x"e6",x"dc",x"c2",x"58"),
   722 => (x"80",x"c1",x"48",x"bf"),
   723 => (x"58",x"ea",x"dc",x"c2"),
   724 => (x"00",x"0c",x"a0",x"27"),
   725 => (x"bf",x"97",x"bf",x"00"),
   726 => (x"c2",x"02",x"9d",x"4d"),
   727 => (x"e5",x"c3",x"87",x"e3"),
   728 => (x"dc",x"c2",x"02",x"ad"),
   729 => (x"e0",x"f2",x"c0",x"87"),
   730 => (x"a3",x"cb",x"4b",x"bf"),
   731 => (x"cf",x"4c",x"11",x"49"),
   732 => (x"d2",x"c1",x"05",x"ac"),
   733 => (x"df",x"49",x"75",x"87"),
   734 => (x"cd",x"89",x"c1",x"99"),
   735 => (x"fa",x"e4",x"c2",x"91"),
   736 => (x"4a",x"a3",x"c1",x"81"),
   737 => (x"a3",x"c3",x"51",x"12"),
   738 => (x"c5",x"51",x"12",x"4a"),
   739 => (x"51",x"12",x"4a",x"a3"),
   740 => (x"12",x"4a",x"a3",x"c7"),
   741 => (x"4a",x"a3",x"c9",x"51"),
   742 => (x"a3",x"ce",x"51",x"12"),
   743 => (x"d0",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"d2"),
   746 => (x"4a",x"a3",x"d4",x"51"),
   747 => (x"a3",x"d6",x"51",x"12"),
   748 => (x"d8",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"dc"),
   751 => (x"4a",x"a3",x"de",x"51"),
   752 => (x"7e",x"c1",x"51",x"12"),
   753 => (x"74",x"87",x"fa",x"c0"),
   754 => (x"05",x"99",x"c8",x"49"),
   755 => (x"74",x"87",x"eb",x"c0"),
   756 => (x"05",x"99",x"d0",x"49"),
   757 => (x"66",x"dc",x"87",x"d1"),
   758 => (x"87",x"cb",x"c0",x"02"),
   759 => (x"66",x"dc",x"49",x"73"),
   760 => (x"02",x"98",x"70",x"0f"),
   761 => (x"6e",x"87",x"d3",x"c0"),
   762 => (x"87",x"c6",x"c0",x"05"),
   763 => (x"48",x"fa",x"e4",x"c2"),
   764 => (x"f2",x"c0",x"50",x"c0"),
   765 => (x"c2",x"48",x"bf",x"e0"),
   766 => (x"e5",x"c2",x"87",x"e1"),
   767 => (x"50",x"c0",x"48",x"c7"),
   768 => (x"f6",x"e4",x"c2",x"7e"),
   769 => (x"dc",x"c2",x"49",x"bf"),
   770 => (x"71",x"4a",x"bf",x"e6"),
   771 => (x"f7",x"fb",x"04",x"aa"),
   772 => (x"d7",x"e9",x"c2",x"87"),
   773 => (x"c8",x"c0",x"05",x"bf"),
   774 => (x"f2",x"e4",x"c2",x"87"),
   775 => (x"f8",x"c1",x"02",x"bf"),
   776 => (x"e2",x"dc",x"c2",x"87"),
   777 => (x"e5",x"ed",x"49",x"bf"),
   778 => (x"c2",x"49",x"70",x"87"),
   779 => (x"c4",x"59",x"e6",x"dc"),
   780 => (x"dc",x"c2",x"48",x"a6"),
   781 => (x"c2",x"78",x"bf",x"e2"),
   782 => (x"02",x"bf",x"f2",x"e4"),
   783 => (x"c4",x"87",x"d8",x"c0"),
   784 => (x"ff",x"cf",x"49",x"66"),
   785 => (x"99",x"f8",x"ff",x"ff"),
   786 => (x"c5",x"c0",x"02",x"a9"),
   787 => (x"c0",x"4c",x"c0",x"87"),
   788 => (x"4c",x"c1",x"87",x"e1"),
   789 => (x"c4",x"87",x"dc",x"c0"),
   790 => (x"ff",x"cf",x"49",x"66"),
   791 => (x"02",x"a9",x"99",x"f8"),
   792 => (x"c8",x"87",x"c8",x"c0"),
   793 => (x"78",x"c0",x"48",x"a6"),
   794 => (x"c8",x"87",x"c5",x"c0"),
   795 => (x"78",x"c1",x"48",x"a6"),
   796 => (x"74",x"4c",x"66",x"c8"),
   797 => (x"e0",x"c0",x"05",x"9c"),
   798 => (x"49",x"66",x"c4",x"87"),
   799 => (x"e4",x"c2",x"89",x"c2"),
   800 => (x"91",x"4a",x"bf",x"ea"),
   801 => (x"bf",x"c3",x"e9",x"c2"),
   802 => (x"de",x"dc",x"c2",x"4a"),
   803 => (x"78",x"a1",x"72",x"48"),
   804 => (x"48",x"e6",x"dc",x"c2"),
   805 => (x"df",x"f9",x"78",x"c0"),
   806 => (x"f4",x"48",x"c0",x"87"),
   807 => (x"87",x"e6",x"eb",x"8e"),
   808 => (x"00",x"00",x"00",x"00"),
   809 => (x"ff",x"ff",x"ff",x"ff"),
   810 => (x"00",x"00",x"0c",x"b0"),
   811 => (x"00",x"00",x"0c",x"b9"),
   812 => (x"33",x"54",x"41",x"46"),
   813 => (x"20",x"20",x"20",x"32"),
   814 => (x"54",x"41",x"46",x"00"),
   815 => (x"20",x"20",x"36",x"31"),
   816 => (x"ff",x"1e",x"00",x"20"),
   817 => (x"ff",x"c3",x"48",x"d4"),
   818 => (x"26",x"48",x"68",x"78"),
   819 => (x"d4",x"ff",x"1e",x"4f"),
   820 => (x"78",x"ff",x"c3",x"48"),
   821 => (x"c0",x"48",x"d0",x"ff"),
   822 => (x"d4",x"ff",x"78",x"e1"),
   823 => (x"c2",x"78",x"d4",x"48"),
   824 => (x"ff",x"48",x"db",x"e9"),
   825 => (x"26",x"50",x"bf",x"d4"),
   826 => (x"d0",x"ff",x"1e",x"4f"),
   827 => (x"78",x"e0",x"c0",x"48"),
   828 => (x"ff",x"1e",x"4f",x"26"),
   829 => (x"49",x"70",x"87",x"cc"),
   830 => (x"87",x"c6",x"02",x"99"),
   831 => (x"05",x"a9",x"fb",x"c0"),
   832 => (x"48",x"71",x"87",x"f1"),
   833 => (x"5e",x"0e",x"4f",x"26"),
   834 => (x"71",x"0e",x"5c",x"5b"),
   835 => (x"fe",x"4c",x"c0",x"4b"),
   836 => (x"49",x"70",x"87",x"f0"),
   837 => (x"f9",x"c0",x"02",x"99"),
   838 => (x"a9",x"ec",x"c0",x"87"),
   839 => (x"87",x"f2",x"c0",x"02"),
   840 => (x"02",x"a9",x"fb",x"c0"),
   841 => (x"cc",x"87",x"eb",x"c0"),
   842 => (x"03",x"ac",x"b7",x"66"),
   843 => (x"66",x"d0",x"87",x"c7"),
   844 => (x"71",x"87",x"c2",x"02"),
   845 => (x"02",x"99",x"71",x"53"),
   846 => (x"84",x"c1",x"87",x"c2"),
   847 => (x"70",x"87",x"c3",x"fe"),
   848 => (x"cd",x"02",x"99",x"49"),
   849 => (x"a9",x"ec",x"c0",x"87"),
   850 => (x"c0",x"87",x"c7",x"02"),
   851 => (x"ff",x"05",x"a9",x"fb"),
   852 => (x"66",x"d0",x"87",x"d5"),
   853 => (x"c0",x"87",x"c3",x"02"),
   854 => (x"ec",x"c0",x"7b",x"97"),
   855 => (x"87",x"c4",x"05",x"a9"),
   856 => (x"87",x"c5",x"4a",x"74"),
   857 => (x"0a",x"c0",x"4a",x"74"),
   858 => (x"c2",x"48",x"72",x"8a"),
   859 => (x"26",x"4d",x"26",x"87"),
   860 => (x"26",x"4b",x"26",x"4c"),
   861 => (x"c9",x"fd",x"1e",x"4f"),
   862 => (x"4a",x"49",x"70",x"87"),
   863 => (x"04",x"aa",x"f0",x"c0"),
   864 => (x"f9",x"c0",x"87",x"c9"),
   865 => (x"87",x"c3",x"01",x"aa"),
   866 => (x"c1",x"8a",x"f0",x"c0"),
   867 => (x"c9",x"04",x"aa",x"c1"),
   868 => (x"aa",x"da",x"c1",x"87"),
   869 => (x"c0",x"87",x"c3",x"01"),
   870 => (x"48",x"72",x"8a",x"f7"),
   871 => (x"5e",x"0e",x"4f",x"26"),
   872 => (x"71",x"0e",x"5c",x"5b"),
   873 => (x"4b",x"d4",x"ff",x"4a"),
   874 => (x"e7",x"c0",x"49",x"72"),
   875 => (x"9c",x"4c",x"70",x"87"),
   876 => (x"c1",x"87",x"c2",x"02"),
   877 => (x"48",x"d0",x"ff",x"8c"),
   878 => (x"d5",x"c1",x"78",x"c5"),
   879 => (x"c6",x"49",x"74",x"7b"),
   880 => (x"d2",x"e4",x"c1",x"31"),
   881 => (x"48",x"4a",x"bf",x"97"),
   882 => (x"7b",x"70",x"b0",x"71"),
   883 => (x"c4",x"48",x"d0",x"ff"),
   884 => (x"87",x"db",x"fe",x"78"),
   885 => (x"5c",x"5b",x"5e",x"0e"),
   886 => (x"86",x"f8",x"0e",x"5d"),
   887 => (x"7e",x"c0",x"4c",x"71"),
   888 => (x"c0",x"87",x"ea",x"fb"),
   889 => (x"c1",x"fa",x"c0",x"4b"),
   890 => (x"c0",x"49",x"bf",x"97"),
   891 => (x"87",x"cf",x"04",x"a9"),
   892 => (x"c1",x"87",x"ff",x"fb"),
   893 => (x"c1",x"fa",x"c0",x"83"),
   894 => (x"ab",x"49",x"bf",x"97"),
   895 => (x"c0",x"87",x"f1",x"06"),
   896 => (x"bf",x"97",x"c1",x"fa"),
   897 => (x"fa",x"87",x"cf",x"02"),
   898 => (x"49",x"70",x"87",x"f8"),
   899 => (x"87",x"c6",x"02",x"99"),
   900 => (x"05",x"a9",x"ec",x"c0"),
   901 => (x"4b",x"c0",x"87",x"f1"),
   902 => (x"70",x"87",x"e7",x"fa"),
   903 => (x"87",x"e2",x"fa",x"4d"),
   904 => (x"fa",x"58",x"a6",x"c8"),
   905 => (x"4a",x"70",x"87",x"dc"),
   906 => (x"a4",x"c8",x"83",x"c1"),
   907 => (x"49",x"69",x"97",x"49"),
   908 => (x"87",x"c7",x"02",x"ad"),
   909 => (x"05",x"ad",x"ff",x"c0"),
   910 => (x"c9",x"87",x"e7",x"c0"),
   911 => (x"69",x"97",x"49",x"a4"),
   912 => (x"a9",x"66",x"c4",x"49"),
   913 => (x"48",x"87",x"c7",x"02"),
   914 => (x"05",x"a8",x"ff",x"c0"),
   915 => (x"a4",x"ca",x"87",x"d4"),
   916 => (x"49",x"69",x"97",x"49"),
   917 => (x"87",x"c6",x"02",x"aa"),
   918 => (x"05",x"aa",x"ff",x"c0"),
   919 => (x"7e",x"c1",x"87",x"c4"),
   920 => (x"ec",x"c0",x"87",x"d0"),
   921 => (x"87",x"c6",x"02",x"ad"),
   922 => (x"05",x"ad",x"fb",x"c0"),
   923 => (x"4b",x"c0",x"87",x"c4"),
   924 => (x"02",x"6e",x"7e",x"c1"),
   925 => (x"f9",x"87",x"e1",x"fe"),
   926 => (x"48",x"73",x"87",x"ef"),
   927 => (x"ec",x"fb",x"8e",x"f8"),
   928 => (x"5e",x"0e",x"00",x"87"),
   929 => (x"0e",x"5d",x"5c",x"5b"),
   930 => (x"4d",x"71",x"86",x"f8"),
   931 => (x"75",x"4b",x"d4",x"ff"),
   932 => (x"e0",x"e9",x"c2",x"1e"),
   933 => (x"87",x"e8",x"e5",x"49"),
   934 => (x"98",x"70",x"86",x"c4"),
   935 => (x"87",x"cc",x"c4",x"02"),
   936 => (x"c1",x"48",x"a6",x"c4"),
   937 => (x"78",x"bf",x"d4",x"e4"),
   938 => (x"f1",x"fb",x"49",x"75"),
   939 => (x"48",x"d0",x"ff",x"87"),
   940 => (x"d6",x"c1",x"78",x"c5"),
   941 => (x"75",x"4a",x"c0",x"7b"),
   942 => (x"7b",x"11",x"49",x"a2"),
   943 => (x"b7",x"cb",x"82",x"c1"),
   944 => (x"87",x"f3",x"04",x"aa"),
   945 => (x"ff",x"c3",x"4a",x"cc"),
   946 => (x"c0",x"82",x"c1",x"7b"),
   947 => (x"04",x"aa",x"b7",x"e0"),
   948 => (x"d0",x"ff",x"87",x"f4"),
   949 => (x"c3",x"78",x"c4",x"48"),
   950 => (x"78",x"c5",x"7b",x"ff"),
   951 => (x"c1",x"7b",x"d3",x"c1"),
   952 => (x"66",x"78",x"c4",x"7b"),
   953 => (x"a8",x"b7",x"c0",x"48"),
   954 => (x"87",x"f0",x"c2",x"06"),
   955 => (x"bf",x"e8",x"e9",x"c2"),
   956 => (x"48",x"66",x"c4",x"4c"),
   957 => (x"a6",x"c8",x"88",x"74"),
   958 => (x"02",x"9c",x"74",x"58"),
   959 => (x"c2",x"87",x"f9",x"c1"),
   960 => (x"c8",x"7e",x"ea",x"dc"),
   961 => (x"c0",x"8c",x"4d",x"c0"),
   962 => (x"c6",x"03",x"ac",x"b7"),
   963 => (x"a4",x"c0",x"c8",x"87"),
   964 => (x"c2",x"4c",x"c0",x"4d"),
   965 => (x"bf",x"97",x"db",x"e9"),
   966 => (x"02",x"99",x"d0",x"49"),
   967 => (x"1e",x"c0",x"87",x"d1"),
   968 => (x"49",x"e0",x"e9",x"c2"),
   969 => (x"c4",x"87",x"cc",x"e8"),
   970 => (x"4a",x"49",x"70",x"86"),
   971 => (x"c2",x"87",x"ee",x"c0"),
   972 => (x"c2",x"1e",x"ea",x"dc"),
   973 => (x"e7",x"49",x"e0",x"e9"),
   974 => (x"86",x"c4",x"87",x"f9"),
   975 => (x"ff",x"4a",x"49",x"70"),
   976 => (x"c5",x"c8",x"48",x"d0"),
   977 => (x"7b",x"d4",x"c1",x"78"),
   978 => (x"7b",x"bf",x"97",x"6e"),
   979 => (x"80",x"c1",x"48",x"6e"),
   980 => (x"8d",x"c1",x"7e",x"70"),
   981 => (x"87",x"f0",x"ff",x"05"),
   982 => (x"c4",x"48",x"d0",x"ff"),
   983 => (x"05",x"9a",x"72",x"78"),
   984 => (x"48",x"c0",x"87",x"c5"),
   985 => (x"c1",x"87",x"c7",x"c1"),
   986 => (x"e0",x"e9",x"c2",x"1e"),
   987 => (x"87",x"e9",x"e5",x"49"),
   988 => (x"9c",x"74",x"86",x"c4"),
   989 => (x"87",x"c7",x"fe",x"05"),
   990 => (x"c0",x"48",x"66",x"c4"),
   991 => (x"d1",x"06",x"a8",x"b7"),
   992 => (x"e0",x"e9",x"c2",x"87"),
   993 => (x"d0",x"78",x"c0",x"48"),
   994 => (x"f4",x"78",x"c0",x"80"),
   995 => (x"ec",x"e9",x"c2",x"80"),
   996 => (x"66",x"c4",x"78",x"bf"),
   997 => (x"a8",x"b7",x"c0",x"48"),
   998 => (x"87",x"d0",x"fd",x"01"),
   999 => (x"c5",x"48",x"d0",x"ff"),
  1000 => (x"7b",x"d3",x"c1",x"78"),
  1001 => (x"78",x"c4",x"7b",x"c0"),
  1002 => (x"87",x"c2",x"48",x"c1"),
  1003 => (x"8e",x"f8",x"48",x"c0"),
  1004 => (x"4c",x"26",x"4d",x"26"),
  1005 => (x"4f",x"26",x"4b",x"26"),
  1006 => (x"5c",x"5b",x"5e",x"0e"),
  1007 => (x"71",x"1e",x"0e",x"5d"),
  1008 => (x"4d",x"4c",x"c0",x"4b"),
  1009 => (x"e8",x"c0",x"04",x"ab"),
  1010 => (x"d4",x"f7",x"c0",x"87"),
  1011 => (x"02",x"9d",x"75",x"1e"),
  1012 => (x"4a",x"c0",x"87",x"c4"),
  1013 => (x"4a",x"c1",x"87",x"c2"),
  1014 => (x"ec",x"eb",x"49",x"72"),
  1015 => (x"70",x"86",x"c4",x"87"),
  1016 => (x"6e",x"84",x"c1",x"7e"),
  1017 => (x"73",x"87",x"c2",x"05"),
  1018 => (x"73",x"85",x"c1",x"4c"),
  1019 => (x"d8",x"ff",x"06",x"ac"),
  1020 => (x"26",x"48",x"6e",x"87"),
  1021 => (x"0e",x"87",x"f9",x"fe"),
  1022 => (x"0e",x"5c",x"5b",x"5e"),
  1023 => (x"66",x"cc",x"4b",x"71"),
  1024 => (x"4c",x"87",x"d8",x"02"),
  1025 => (x"02",x"8c",x"f0",x"c0"),
  1026 => (x"4a",x"74",x"87",x"d8"),
  1027 => (x"d1",x"02",x"8a",x"c1"),
  1028 => (x"cd",x"02",x"8a",x"87"),
  1029 => (x"c9",x"02",x"8a",x"87"),
  1030 => (x"73",x"87",x"d9",x"87"),
  1031 => (x"87",x"e2",x"f9",x"49"),
  1032 => (x"1e",x"74",x"87",x"d2"),
  1033 => (x"d7",x"c1",x"49",x"c0"),
  1034 => (x"1e",x"74",x"87",x"f5"),
  1035 => (x"d7",x"c1",x"49",x"73"),
  1036 => (x"86",x"c8",x"87",x"ed"),
  1037 => (x"0e",x"87",x"fb",x"fd"),
  1038 => (x"5d",x"5c",x"5b",x"5e"),
  1039 => (x"4c",x"71",x"1e",x"0e"),
  1040 => (x"c2",x"91",x"de",x"49"),
  1041 => (x"71",x"4d",x"c8",x"ea"),
  1042 => (x"02",x"6d",x"97",x"85"),
  1043 => (x"c2",x"87",x"dd",x"c1"),
  1044 => (x"4a",x"bf",x"f4",x"e9"),
  1045 => (x"49",x"72",x"82",x"74"),
  1046 => (x"70",x"87",x"dd",x"fd"),
  1047 => (x"02",x"98",x"48",x"7e"),
  1048 => (x"c2",x"87",x"f2",x"c0"),
  1049 => (x"70",x"4b",x"fc",x"e9"),
  1050 => (x"ff",x"49",x"cb",x"4a"),
  1051 => (x"74",x"87",x"f8",x"c0"),
  1052 => (x"c1",x"93",x"cb",x"4b"),
  1053 => (x"c4",x"83",x"e6",x"e4"),
  1054 => (x"f0",x"c2",x"c1",x"83"),
  1055 => (x"c1",x"49",x"74",x"7b"),
  1056 => (x"75",x"87",x"d3",x"c0"),
  1057 => (x"d3",x"e4",x"c1",x"7b"),
  1058 => (x"1e",x"49",x"bf",x"97"),
  1059 => (x"49",x"fc",x"e9",x"c2"),
  1060 => (x"c4",x"87",x"e4",x"fd"),
  1061 => (x"c0",x"49",x"74",x"86"),
  1062 => (x"c0",x"87",x"fb",x"ff"),
  1063 => (x"da",x"c1",x"c1",x"49"),
  1064 => (x"dc",x"e9",x"c2",x"87"),
  1065 => (x"c1",x"78",x"c0",x"48"),
  1066 => (x"87",x"de",x"de",x"49"),
  1067 => (x"87",x"c0",x"fc",x"26"),
  1068 => (x"64",x"61",x"6f",x"4c"),
  1069 => (x"2e",x"67",x"6e",x"69"),
  1070 => (x"0e",x"00",x"2e",x"2e"),
  1071 => (x"0e",x"5c",x"5b",x"5e"),
  1072 => (x"c2",x"4a",x"4b",x"71"),
  1073 => (x"82",x"bf",x"f4",x"e9"),
  1074 => (x"eb",x"fb",x"49",x"72"),
  1075 => (x"9c",x"4c",x"70",x"87"),
  1076 => (x"49",x"87",x"c4",x"02"),
  1077 => (x"c2",x"87",x"fa",x"e6"),
  1078 => (x"c0",x"48",x"f4",x"e9"),
  1079 => (x"dd",x"49",x"c1",x"78"),
  1080 => (x"cd",x"fb",x"87",x"e8"),
  1081 => (x"5b",x"5e",x"0e",x"87"),
  1082 => (x"f4",x"0e",x"5d",x"5c"),
  1083 => (x"ea",x"dc",x"c2",x"86"),
  1084 => (x"c4",x"4c",x"c0",x"4d"),
  1085 => (x"78",x"c0",x"48",x"a6"),
  1086 => (x"bf",x"f4",x"e9",x"c2"),
  1087 => (x"06",x"a9",x"c0",x"49"),
  1088 => (x"c2",x"87",x"c1",x"c1"),
  1089 => (x"98",x"48",x"ea",x"dc"),
  1090 => (x"87",x"f8",x"c0",x"02"),
  1091 => (x"1e",x"d4",x"f7",x"c0"),
  1092 => (x"c7",x"02",x"66",x"c8"),
  1093 => (x"48",x"a6",x"c4",x"87"),
  1094 => (x"87",x"c5",x"78",x"c0"),
  1095 => (x"c1",x"48",x"a6",x"c4"),
  1096 => (x"49",x"66",x"c4",x"78"),
  1097 => (x"c4",x"87",x"e2",x"e6"),
  1098 => (x"c1",x"4d",x"70",x"86"),
  1099 => (x"48",x"66",x"c4",x"84"),
  1100 => (x"a6",x"c8",x"80",x"c1"),
  1101 => (x"f4",x"e9",x"c2",x"58"),
  1102 => (x"03",x"ac",x"49",x"bf"),
  1103 => (x"9d",x"75",x"87",x"c6"),
  1104 => (x"87",x"c8",x"ff",x"05"),
  1105 => (x"9d",x"75",x"4c",x"c0"),
  1106 => (x"87",x"e0",x"c3",x"02"),
  1107 => (x"1e",x"d4",x"f7",x"c0"),
  1108 => (x"c7",x"02",x"66",x"c8"),
  1109 => (x"48",x"a6",x"cc",x"87"),
  1110 => (x"87",x"c5",x"78",x"c0"),
  1111 => (x"c1",x"48",x"a6",x"cc"),
  1112 => (x"49",x"66",x"cc",x"78"),
  1113 => (x"c4",x"87",x"e2",x"e5"),
  1114 => (x"48",x"7e",x"70",x"86"),
  1115 => (x"e8",x"c2",x"02",x"98"),
  1116 => (x"81",x"cb",x"49",x"87"),
  1117 => (x"d0",x"49",x"69",x"97"),
  1118 => (x"d6",x"c1",x"02",x"99"),
  1119 => (x"fb",x"c2",x"c1",x"87"),
  1120 => (x"cb",x"49",x"74",x"4a"),
  1121 => (x"e6",x"e4",x"c1",x"91"),
  1122 => (x"c8",x"79",x"72",x"81"),
  1123 => (x"51",x"ff",x"c3",x"81"),
  1124 => (x"91",x"de",x"49",x"74"),
  1125 => (x"4d",x"c8",x"ea",x"c2"),
  1126 => (x"c1",x"c2",x"85",x"71"),
  1127 => (x"a5",x"c1",x"7d",x"97"),
  1128 => (x"51",x"e0",x"c0",x"49"),
  1129 => (x"97",x"fa",x"e4",x"c2"),
  1130 => (x"87",x"d2",x"02",x"bf"),
  1131 => (x"a5",x"c2",x"84",x"c1"),
  1132 => (x"fa",x"e4",x"c2",x"4b"),
  1133 => (x"fe",x"49",x"db",x"4a"),
  1134 => (x"c1",x"87",x"ec",x"fb"),
  1135 => (x"a5",x"cd",x"87",x"db"),
  1136 => (x"c1",x"51",x"c0",x"49"),
  1137 => (x"4b",x"a5",x"c2",x"84"),
  1138 => (x"49",x"cb",x"4a",x"6e"),
  1139 => (x"87",x"d7",x"fb",x"fe"),
  1140 => (x"c1",x"87",x"c6",x"c1"),
  1141 => (x"74",x"4a",x"f7",x"c0"),
  1142 => (x"c1",x"91",x"cb",x"49"),
  1143 => (x"72",x"81",x"e6",x"e4"),
  1144 => (x"fa",x"e4",x"c2",x"79"),
  1145 => (x"d8",x"02",x"bf",x"97"),
  1146 => (x"de",x"49",x"74",x"87"),
  1147 => (x"c2",x"84",x"c1",x"91"),
  1148 => (x"71",x"4b",x"c8",x"ea"),
  1149 => (x"fa",x"e4",x"c2",x"83"),
  1150 => (x"fe",x"49",x"dd",x"4a"),
  1151 => (x"d8",x"87",x"e8",x"fa"),
  1152 => (x"de",x"4b",x"74",x"87"),
  1153 => (x"c8",x"ea",x"c2",x"93"),
  1154 => (x"49",x"a3",x"cb",x"83"),
  1155 => (x"84",x"c1",x"51",x"c0"),
  1156 => (x"cb",x"4a",x"6e",x"73"),
  1157 => (x"ce",x"fa",x"fe",x"49"),
  1158 => (x"48",x"66",x"c4",x"87"),
  1159 => (x"a6",x"c8",x"80",x"c1"),
  1160 => (x"03",x"ac",x"c7",x"58"),
  1161 => (x"6e",x"87",x"c5",x"c0"),
  1162 => (x"87",x"e0",x"fc",x"05"),
  1163 => (x"8e",x"f4",x"48",x"74"),
  1164 => (x"1e",x"87",x"fd",x"f5"),
  1165 => (x"4b",x"71",x"1e",x"73"),
  1166 => (x"c1",x"91",x"cb",x"49"),
  1167 => (x"c8",x"81",x"e6",x"e4"),
  1168 => (x"e4",x"c1",x"4a",x"a1"),
  1169 => (x"50",x"12",x"48",x"d2"),
  1170 => (x"c0",x"4a",x"a1",x"c9"),
  1171 => (x"12",x"48",x"c1",x"fa"),
  1172 => (x"c1",x"81",x"ca",x"50"),
  1173 => (x"11",x"48",x"d3",x"e4"),
  1174 => (x"d3",x"e4",x"c1",x"50"),
  1175 => (x"1e",x"49",x"bf",x"97"),
  1176 => (x"d2",x"f6",x"49",x"c0"),
  1177 => (x"dc",x"e9",x"c2",x"87"),
  1178 => (x"c1",x"78",x"de",x"48"),
  1179 => (x"87",x"da",x"d7",x"49"),
  1180 => (x"87",x"c0",x"f5",x"26"),
  1181 => (x"49",x"4a",x"71",x"1e"),
  1182 => (x"e4",x"c1",x"91",x"cb"),
  1183 => (x"81",x"c8",x"81",x"e6"),
  1184 => (x"e9",x"c2",x"48",x"11"),
  1185 => (x"e9",x"c2",x"58",x"e0"),
  1186 => (x"78",x"c0",x"48",x"f4"),
  1187 => (x"f9",x"d6",x"49",x"c1"),
  1188 => (x"1e",x"4f",x"26",x"87"),
  1189 => (x"f9",x"c0",x"49",x"c0"),
  1190 => (x"4f",x"26",x"87",x"e1"),
  1191 => (x"02",x"99",x"71",x"1e"),
  1192 => (x"e5",x"c1",x"87",x"d2"),
  1193 => (x"50",x"c0",x"48",x"fb"),
  1194 => (x"c9",x"c1",x"80",x"f7"),
  1195 => (x"e4",x"c1",x"40",x"f4"),
  1196 => (x"87",x"ce",x"78",x"df"),
  1197 => (x"48",x"f7",x"e5",x"c1"),
  1198 => (x"78",x"d8",x"e4",x"c1"),
  1199 => (x"ca",x"c1",x"80",x"fc"),
  1200 => (x"4f",x"26",x"78",x"d3"),
  1201 => (x"5c",x"5b",x"5e",x"0e"),
  1202 => (x"86",x"f4",x"0e",x"5d"),
  1203 => (x"cb",x"49",x"4d",x"71"),
  1204 => (x"e6",x"e4",x"c1",x"91"),
  1205 => (x"4a",x"a1",x"c8",x"81"),
  1206 => (x"c4",x"7e",x"a1",x"ca"),
  1207 => (x"ed",x"c2",x"48",x"a6"),
  1208 => (x"6e",x"78",x"bf",x"e4"),
  1209 => (x"c4",x"4b",x"bf",x"97"),
  1210 => (x"28",x"73",x"48",x"66"),
  1211 => (x"12",x"4c",x"4b",x"70"),
  1212 => (x"58",x"a6",x"cc",x"48"),
  1213 => (x"84",x"c1",x"9c",x"70"),
  1214 => (x"69",x"97",x"81",x"c9"),
  1215 => (x"04",x"ac",x"b7",x"49"),
  1216 => (x"4c",x"c0",x"87",x"c2"),
  1217 => (x"4a",x"bf",x"97",x"6e"),
  1218 => (x"72",x"49",x"66",x"c8"),
  1219 => (x"c4",x"b9",x"ff",x"31"),
  1220 => (x"48",x"74",x"99",x"66"),
  1221 => (x"4a",x"70",x"30",x"72"),
  1222 => (x"c2",x"b0",x"71",x"48"),
  1223 => (x"c0",x"58",x"e8",x"ed"),
  1224 => (x"c0",x"87",x"f3",x"e3"),
  1225 => (x"87",x"e2",x"d4",x"49"),
  1226 => (x"f5",x"c0",x"49",x"75"),
  1227 => (x"8e",x"f4",x"87",x"e8"),
  1228 => (x"1e",x"87",x"fd",x"f1"),
  1229 => (x"4b",x"71",x"1e",x"73"),
  1230 => (x"87",x"c8",x"fe",x"49"),
  1231 => (x"c3",x"fe",x"49",x"73"),
  1232 => (x"87",x"f0",x"f1",x"87"),
  1233 => (x"71",x"1e",x"73",x"1e"),
  1234 => (x"4a",x"a3",x"c6",x"4b"),
  1235 => (x"c1",x"87",x"db",x"02"),
  1236 => (x"87",x"d6",x"02",x"8a"),
  1237 => (x"da",x"c1",x"02",x"8a"),
  1238 => (x"c0",x"02",x"8a",x"87"),
  1239 => (x"02",x"8a",x"87",x"fc"),
  1240 => (x"8a",x"87",x"e1",x"c0"),
  1241 => (x"c1",x"87",x"cb",x"02"),
  1242 => (x"49",x"c7",x"87",x"db"),
  1243 => (x"c1",x"87",x"c5",x"fc"),
  1244 => (x"e9",x"c2",x"87",x"de"),
  1245 => (x"c1",x"02",x"bf",x"f4"),
  1246 => (x"c1",x"48",x"87",x"cb"),
  1247 => (x"f8",x"e9",x"c2",x"88"),
  1248 => (x"87",x"c1",x"c1",x"58"),
  1249 => (x"bf",x"f8",x"e9",x"c2"),
  1250 => (x"87",x"f9",x"c0",x"02"),
  1251 => (x"bf",x"f4",x"e9",x"c2"),
  1252 => (x"c2",x"80",x"c1",x"48"),
  1253 => (x"c0",x"58",x"f8",x"e9"),
  1254 => (x"e9",x"c2",x"87",x"eb"),
  1255 => (x"c6",x"49",x"bf",x"f4"),
  1256 => (x"f8",x"e9",x"c2",x"89"),
  1257 => (x"a9",x"b7",x"c0",x"59"),
  1258 => (x"c2",x"87",x"da",x"03"),
  1259 => (x"c0",x"48",x"f4",x"e9"),
  1260 => (x"c2",x"87",x"d2",x"78"),
  1261 => (x"02",x"bf",x"f8",x"e9"),
  1262 => (x"e9",x"c2",x"87",x"cb"),
  1263 => (x"c6",x"48",x"bf",x"f4"),
  1264 => (x"f8",x"e9",x"c2",x"80"),
  1265 => (x"d2",x"49",x"c0",x"58"),
  1266 => (x"49",x"73",x"87",x"c0"),
  1267 => (x"87",x"c6",x"f3",x"c0"),
  1268 => (x"0e",x"87",x"e1",x"ef"),
  1269 => (x"5d",x"5c",x"5b",x"5e"),
  1270 => (x"86",x"d0",x"ff",x"0e"),
  1271 => (x"c8",x"59",x"a6",x"dc"),
  1272 => (x"78",x"c0",x"48",x"a6"),
  1273 => (x"c4",x"c1",x"80",x"c4"),
  1274 => (x"80",x"c4",x"78",x"66"),
  1275 => (x"80",x"c4",x"78",x"c1"),
  1276 => (x"e9",x"c2",x"78",x"c1"),
  1277 => (x"78",x"c1",x"48",x"f8"),
  1278 => (x"bf",x"dc",x"e9",x"c2"),
  1279 => (x"05",x"a8",x"de",x"48"),
  1280 => (x"e0",x"f3",x"87",x"cb"),
  1281 => (x"cc",x"49",x"70",x"87"),
  1282 => (x"fc",x"cf",x"59",x"a6"),
  1283 => (x"87",x"fd",x"e2",x"87"),
  1284 => (x"e2",x"87",x"df",x"e3"),
  1285 => (x"4c",x"70",x"87",x"ec"),
  1286 => (x"02",x"ac",x"fb",x"c0"),
  1287 => (x"d8",x"87",x"fb",x"c1"),
  1288 => (x"ed",x"c1",x"05",x"66"),
  1289 => (x"66",x"c0",x"c1",x"87"),
  1290 => (x"6a",x"82",x"c4",x"4a"),
  1291 => (x"c1",x"1e",x"72",x"7e"),
  1292 => (x"c4",x"48",x"fe",x"e0"),
  1293 => (x"a1",x"c8",x"49",x"66"),
  1294 => (x"71",x"41",x"20",x"4a"),
  1295 => (x"87",x"f9",x"05",x"aa"),
  1296 => (x"4a",x"26",x"51",x"10"),
  1297 => (x"48",x"66",x"c0",x"c1"),
  1298 => (x"78",x"f3",x"c8",x"c1"),
  1299 => (x"81",x"c7",x"49",x"6a"),
  1300 => (x"c0",x"c1",x"51",x"74"),
  1301 => (x"81",x"c8",x"49",x"66"),
  1302 => (x"c0",x"c1",x"51",x"c1"),
  1303 => (x"81",x"c9",x"49",x"66"),
  1304 => (x"c0",x"c1",x"51",x"c0"),
  1305 => (x"81",x"ca",x"49",x"66"),
  1306 => (x"1e",x"c1",x"51",x"c0"),
  1307 => (x"49",x"6a",x"1e",x"d8"),
  1308 => (x"d1",x"e2",x"81",x"c8"),
  1309 => (x"c1",x"86",x"c8",x"87"),
  1310 => (x"c0",x"48",x"66",x"c4"),
  1311 => (x"87",x"c7",x"01",x"a8"),
  1312 => (x"c1",x"48",x"a6",x"c8"),
  1313 => (x"c1",x"87",x"ce",x"78"),
  1314 => (x"c1",x"48",x"66",x"c4"),
  1315 => (x"58",x"a6",x"d0",x"88"),
  1316 => (x"dd",x"e1",x"87",x"c3"),
  1317 => (x"48",x"a6",x"d0",x"87"),
  1318 => (x"9c",x"74",x"78",x"c2"),
  1319 => (x"87",x"e5",x"cd",x"02"),
  1320 => (x"c1",x"48",x"66",x"c8"),
  1321 => (x"03",x"a8",x"66",x"c8"),
  1322 => (x"dc",x"87",x"da",x"cd"),
  1323 => (x"78",x"c0",x"48",x"a6"),
  1324 => (x"78",x"c0",x"80",x"e8"),
  1325 => (x"70",x"87",x"cb",x"e0"),
  1326 => (x"ac",x"d0",x"c1",x"4c"),
  1327 => (x"87",x"da",x"c2",x"05"),
  1328 => (x"e2",x"7e",x"66",x"c4"),
  1329 => (x"49",x"70",x"87",x"ef"),
  1330 => (x"ff",x"59",x"a6",x"c8"),
  1331 => (x"70",x"87",x"f3",x"df"),
  1332 => (x"ac",x"ec",x"c0",x"4c"),
  1333 => (x"87",x"ed",x"c1",x"05"),
  1334 => (x"cb",x"49",x"66",x"c8"),
  1335 => (x"66",x"c0",x"c1",x"91"),
  1336 => (x"4a",x"a1",x"c4",x"81"),
  1337 => (x"a1",x"c8",x"4d",x"6a"),
  1338 => (x"52",x"66",x"c4",x"4a"),
  1339 => (x"79",x"f4",x"c9",x"c1"),
  1340 => (x"87",x"ce",x"df",x"ff"),
  1341 => (x"02",x"9c",x"4c",x"70"),
  1342 => (x"fb",x"c0",x"87",x"d9"),
  1343 => (x"87",x"d3",x"02",x"ac"),
  1344 => (x"de",x"ff",x"55",x"74"),
  1345 => (x"4c",x"70",x"87",x"fc"),
  1346 => (x"87",x"c7",x"02",x"9c"),
  1347 => (x"05",x"ac",x"fb",x"c0"),
  1348 => (x"c0",x"87",x"ed",x"ff"),
  1349 => (x"c1",x"c2",x"55",x"e0"),
  1350 => (x"7d",x"97",x"c0",x"55"),
  1351 => (x"6e",x"49",x"66",x"d8"),
  1352 => (x"87",x"db",x"05",x"a9"),
  1353 => (x"cc",x"48",x"66",x"c8"),
  1354 => (x"ca",x"04",x"a8",x"66"),
  1355 => (x"48",x"66",x"c8",x"87"),
  1356 => (x"a6",x"cc",x"80",x"c1"),
  1357 => (x"cc",x"87",x"c8",x"58"),
  1358 => (x"88",x"c1",x"48",x"66"),
  1359 => (x"ff",x"58",x"a6",x"d0"),
  1360 => (x"70",x"87",x"ff",x"dd"),
  1361 => (x"ac",x"d0",x"c1",x"4c"),
  1362 => (x"d4",x"87",x"c8",x"05"),
  1363 => (x"80",x"c1",x"48",x"66"),
  1364 => (x"c1",x"58",x"a6",x"d8"),
  1365 => (x"fd",x"02",x"ac",x"d0"),
  1366 => (x"e0",x"c0",x"87",x"e6"),
  1367 => (x"66",x"d8",x"48",x"a6"),
  1368 => (x"48",x"66",x"c4",x"78"),
  1369 => (x"a8",x"66",x"e0",x"c0"),
  1370 => (x"87",x"eb",x"c9",x"05"),
  1371 => (x"48",x"a6",x"e4",x"c0"),
  1372 => (x"48",x"74",x"78",x"c0"),
  1373 => (x"70",x"88",x"fb",x"c0"),
  1374 => (x"02",x"98",x"48",x"7e"),
  1375 => (x"48",x"87",x"ed",x"c9"),
  1376 => (x"7e",x"70",x"88",x"cb"),
  1377 => (x"c1",x"02",x"98",x"48"),
  1378 => (x"c9",x"48",x"87",x"cd"),
  1379 => (x"48",x"7e",x"70",x"88"),
  1380 => (x"c1",x"c4",x"02",x"98"),
  1381 => (x"88",x"c4",x"48",x"87"),
  1382 => (x"98",x"48",x"7e",x"70"),
  1383 => (x"48",x"87",x"ce",x"02"),
  1384 => (x"7e",x"70",x"88",x"c1"),
  1385 => (x"c3",x"02",x"98",x"48"),
  1386 => (x"e1",x"c8",x"87",x"ec"),
  1387 => (x"48",x"a6",x"dc",x"87"),
  1388 => (x"ff",x"78",x"f0",x"c0"),
  1389 => (x"70",x"87",x"cb",x"dc"),
  1390 => (x"ac",x"ec",x"c0",x"4c"),
  1391 => (x"87",x"c4",x"c0",x"02"),
  1392 => (x"5c",x"a6",x"e0",x"c0"),
  1393 => (x"02",x"ac",x"ec",x"c0"),
  1394 => (x"db",x"ff",x"87",x"cd"),
  1395 => (x"4c",x"70",x"87",x"f4"),
  1396 => (x"05",x"ac",x"ec",x"c0"),
  1397 => (x"c0",x"87",x"f3",x"ff"),
  1398 => (x"c0",x"02",x"ac",x"ec"),
  1399 => (x"db",x"ff",x"87",x"c4"),
  1400 => (x"1e",x"c0",x"87",x"e0"),
  1401 => (x"66",x"d0",x"1e",x"ca"),
  1402 => (x"c1",x"91",x"cb",x"49"),
  1403 => (x"71",x"48",x"66",x"c8"),
  1404 => (x"58",x"a6",x"cc",x"80"),
  1405 => (x"c4",x"48",x"66",x"c8"),
  1406 => (x"58",x"a6",x"d0",x"80"),
  1407 => (x"49",x"bf",x"66",x"cc"),
  1408 => (x"87",x"c2",x"dc",x"ff"),
  1409 => (x"1e",x"de",x"1e",x"c1"),
  1410 => (x"49",x"bf",x"66",x"d4"),
  1411 => (x"87",x"f6",x"db",x"ff"),
  1412 => (x"49",x"70",x"86",x"d0"),
  1413 => (x"c0",x"89",x"09",x"c0"),
  1414 => (x"c0",x"59",x"a6",x"ec"),
  1415 => (x"c0",x"48",x"66",x"e8"),
  1416 => (x"ee",x"c0",x"06",x"a8"),
  1417 => (x"66",x"e8",x"c0",x"87"),
  1418 => (x"03",x"a8",x"dd",x"48"),
  1419 => (x"c4",x"87",x"e4",x"c0"),
  1420 => (x"c0",x"49",x"bf",x"66"),
  1421 => (x"c0",x"81",x"66",x"e8"),
  1422 => (x"e8",x"c0",x"51",x"e0"),
  1423 => (x"81",x"c1",x"49",x"66"),
  1424 => (x"81",x"bf",x"66",x"c4"),
  1425 => (x"c0",x"51",x"c1",x"c2"),
  1426 => (x"c2",x"49",x"66",x"e8"),
  1427 => (x"bf",x"66",x"c4",x"81"),
  1428 => (x"6e",x"51",x"c0",x"81"),
  1429 => (x"f3",x"c8",x"c1",x"48"),
  1430 => (x"c8",x"49",x"6e",x"78"),
  1431 => (x"51",x"66",x"d0",x"81"),
  1432 => (x"81",x"c9",x"49",x"6e"),
  1433 => (x"6e",x"51",x"66",x"d4"),
  1434 => (x"dc",x"81",x"ca",x"49"),
  1435 => (x"66",x"d0",x"51",x"66"),
  1436 => (x"d4",x"80",x"c1",x"48"),
  1437 => (x"66",x"c8",x"58",x"a6"),
  1438 => (x"a8",x"66",x"cc",x"48"),
  1439 => (x"87",x"cb",x"c0",x"04"),
  1440 => (x"c1",x"48",x"66",x"c8"),
  1441 => (x"58",x"a6",x"cc",x"80"),
  1442 => (x"cc",x"87",x"e1",x"c5"),
  1443 => (x"88",x"c1",x"48",x"66"),
  1444 => (x"c5",x"58",x"a6",x"d0"),
  1445 => (x"db",x"ff",x"87",x"d6"),
  1446 => (x"49",x"70",x"87",x"db"),
  1447 => (x"59",x"a6",x"ec",x"c0"),
  1448 => (x"87",x"d1",x"db",x"ff"),
  1449 => (x"e0",x"c0",x"49",x"70"),
  1450 => (x"66",x"dc",x"59",x"a6"),
  1451 => (x"a8",x"ec",x"c0",x"48"),
  1452 => (x"87",x"ca",x"c0",x"05"),
  1453 => (x"c0",x"48",x"a6",x"dc"),
  1454 => (x"c0",x"78",x"66",x"e8"),
  1455 => (x"d8",x"ff",x"87",x"c4"),
  1456 => (x"66",x"c8",x"87",x"c0"),
  1457 => (x"c1",x"91",x"cb",x"49"),
  1458 => (x"71",x"48",x"66",x"c0"),
  1459 => (x"4a",x"7e",x"70",x"80"),
  1460 => (x"49",x"6e",x"82",x"c8"),
  1461 => (x"e8",x"c0",x"81",x"ca"),
  1462 => (x"66",x"dc",x"51",x"66"),
  1463 => (x"c0",x"81",x"c1",x"49"),
  1464 => (x"c1",x"89",x"66",x"e8"),
  1465 => (x"70",x"30",x"71",x"48"),
  1466 => (x"71",x"89",x"c1",x"49"),
  1467 => (x"ed",x"c2",x"7a",x"97"),
  1468 => (x"c0",x"49",x"bf",x"e4"),
  1469 => (x"97",x"29",x"66",x"e8"),
  1470 => (x"71",x"48",x"4a",x"6a"),
  1471 => (x"a6",x"f0",x"c0",x"98"),
  1472 => (x"c4",x"49",x"6e",x"58"),
  1473 => (x"c0",x"4d",x"69",x"81"),
  1474 => (x"c4",x"48",x"66",x"e0"),
  1475 => (x"c0",x"02",x"a8",x"66"),
  1476 => (x"a6",x"c4",x"87",x"c8"),
  1477 => (x"c0",x"78",x"c0",x"48"),
  1478 => (x"a6",x"c4",x"87",x"c5"),
  1479 => (x"c4",x"78",x"c1",x"48"),
  1480 => (x"e0",x"c0",x"1e",x"66"),
  1481 => (x"ff",x"49",x"75",x"1e"),
  1482 => (x"c8",x"87",x"db",x"d7"),
  1483 => (x"c0",x"4c",x"70",x"86"),
  1484 => (x"c1",x"06",x"ac",x"b7"),
  1485 => (x"85",x"74",x"87",x"d4"),
  1486 => (x"74",x"49",x"e0",x"c0"),
  1487 => (x"c1",x"4b",x"75",x"89"),
  1488 => (x"71",x"4a",x"c7",x"e1"),
  1489 => (x"87",x"df",x"e5",x"fe"),
  1490 => (x"e4",x"c0",x"85",x"c2"),
  1491 => (x"80",x"c1",x"48",x"66"),
  1492 => (x"58",x"a6",x"e8",x"c0"),
  1493 => (x"49",x"66",x"ec",x"c0"),
  1494 => (x"a9",x"70",x"81",x"c1"),
  1495 => (x"87",x"c8",x"c0",x"02"),
  1496 => (x"c0",x"48",x"a6",x"c4"),
  1497 => (x"87",x"c5",x"c0",x"78"),
  1498 => (x"c1",x"48",x"a6",x"c4"),
  1499 => (x"1e",x"66",x"c4",x"78"),
  1500 => (x"c0",x"49",x"a4",x"c2"),
  1501 => (x"88",x"71",x"48",x"e0"),
  1502 => (x"75",x"1e",x"49",x"70"),
  1503 => (x"c5",x"d6",x"ff",x"49"),
  1504 => (x"c0",x"86",x"c8",x"87"),
  1505 => (x"ff",x"01",x"a8",x"b7"),
  1506 => (x"e4",x"c0",x"87",x"c0"),
  1507 => (x"d1",x"c0",x"02",x"66"),
  1508 => (x"c9",x"49",x"6e",x"87"),
  1509 => (x"66",x"e4",x"c0",x"81"),
  1510 => (x"c1",x"48",x"6e",x"51"),
  1511 => (x"c0",x"78",x"c4",x"cb"),
  1512 => (x"49",x"6e",x"87",x"cc"),
  1513 => (x"51",x"c2",x"81",x"c9"),
  1514 => (x"cc",x"c1",x"48",x"6e"),
  1515 => (x"66",x"c8",x"78",x"f3"),
  1516 => (x"a8",x"66",x"cc",x"48"),
  1517 => (x"87",x"cb",x"c0",x"04"),
  1518 => (x"c1",x"48",x"66",x"c8"),
  1519 => (x"58",x"a6",x"cc",x"80"),
  1520 => (x"cc",x"87",x"e9",x"c0"),
  1521 => (x"88",x"c1",x"48",x"66"),
  1522 => (x"c0",x"58",x"a6",x"d0"),
  1523 => (x"d4",x"ff",x"87",x"de"),
  1524 => (x"4c",x"70",x"87",x"e0"),
  1525 => (x"c1",x"87",x"d5",x"c0"),
  1526 => (x"c0",x"05",x"ac",x"c6"),
  1527 => (x"66",x"d0",x"87",x"c8"),
  1528 => (x"d4",x"80",x"c1",x"48"),
  1529 => (x"d4",x"ff",x"58",x"a6"),
  1530 => (x"4c",x"70",x"87",x"c8"),
  1531 => (x"c1",x"48",x"66",x"d4"),
  1532 => (x"58",x"a6",x"d8",x"80"),
  1533 => (x"c0",x"02",x"9c",x"74"),
  1534 => (x"66",x"c8",x"87",x"cb"),
  1535 => (x"66",x"c8",x"c1",x"48"),
  1536 => (x"e6",x"f2",x"04",x"a8"),
  1537 => (x"e0",x"d3",x"ff",x"87"),
  1538 => (x"48",x"66",x"c8",x"87"),
  1539 => (x"c0",x"03",x"a8",x"c7"),
  1540 => (x"e9",x"c2",x"87",x"e5"),
  1541 => (x"78",x"c0",x"48",x"f8"),
  1542 => (x"cb",x"49",x"66",x"c8"),
  1543 => (x"66",x"c0",x"c1",x"91"),
  1544 => (x"4a",x"a1",x"c4",x"81"),
  1545 => (x"52",x"c0",x"4a",x"6a"),
  1546 => (x"48",x"66",x"c8",x"79"),
  1547 => (x"a6",x"cc",x"80",x"c1"),
  1548 => (x"04",x"a8",x"c7",x"58"),
  1549 => (x"ff",x"87",x"db",x"ff"),
  1550 => (x"dd",x"ff",x"8e",x"d0"),
  1551 => (x"6f",x"4c",x"87",x"f2"),
  1552 => (x"2a",x"20",x"64",x"61"),
  1553 => (x"3a",x"00",x"20",x"2e"),
  1554 => (x"73",x"1e",x"00",x"20"),
  1555 => (x"9b",x"4b",x"71",x"1e"),
  1556 => (x"c2",x"87",x"c6",x"02"),
  1557 => (x"c0",x"48",x"f4",x"e9"),
  1558 => (x"c2",x"1e",x"c7",x"78"),
  1559 => (x"49",x"bf",x"f4",x"e9"),
  1560 => (x"e6",x"e4",x"c1",x"1e"),
  1561 => (x"dc",x"e9",x"c2",x"1e"),
  1562 => (x"e6",x"ed",x"49",x"bf"),
  1563 => (x"c2",x"86",x"cc",x"87"),
  1564 => (x"49",x"bf",x"dc",x"e9"),
  1565 => (x"73",x"87",x"e5",x"e8"),
  1566 => (x"87",x"c8",x"02",x"9b"),
  1567 => (x"49",x"e6",x"e4",x"c1"),
  1568 => (x"87",x"e4",x"e1",x"c0"),
  1569 => (x"87",x"ec",x"dc",x"ff"),
  1570 => (x"87",x"d4",x"c7",x"1e"),
  1571 => (x"f9",x"fe",x"49",x"c1"),
  1572 => (x"fa",x"e8",x"fe",x"87"),
  1573 => (x"02",x"98",x"70",x"87"),
  1574 => (x"f1",x"fe",x"87",x"cd"),
  1575 => (x"98",x"70",x"87",x"f5"),
  1576 => (x"c1",x"87",x"c4",x"02"),
  1577 => (x"c0",x"87",x"c2",x"4a"),
  1578 => (x"05",x"9a",x"72",x"4a"),
  1579 => (x"1e",x"c0",x"87",x"ce"),
  1580 => (x"49",x"d9",x"e3",x"c1"),
  1581 => (x"87",x"dd",x"ee",x"c0"),
  1582 => (x"87",x"fe",x"86",x"c4"),
  1583 => (x"e3",x"c1",x"1e",x"c0"),
  1584 => (x"ee",x"c0",x"49",x"e4"),
  1585 => (x"1e",x"c0",x"87",x"cf"),
  1586 => (x"87",x"d4",x"f7",x"c0"),
  1587 => (x"ee",x"c0",x"49",x"70"),
  1588 => (x"ca",x"c3",x"87",x"c3"),
  1589 => (x"26",x"8e",x"f8",x"87"),
  1590 => (x"20",x"44",x"53",x"4f"),
  1591 => (x"6c",x"69",x"61",x"66"),
  1592 => (x"00",x"2e",x"64",x"65"),
  1593 => (x"74",x"6f",x"6f",x"42"),
  1594 => (x"2e",x"67",x"6e",x"69"),
  1595 => (x"1e",x"00",x"2e",x"2e"),
  1596 => (x"87",x"f2",x"e4",x"c0"),
  1597 => (x"87",x"d7",x"f1",x"c0"),
  1598 => (x"4f",x"26",x"87",x"f6"),
  1599 => (x"f4",x"e9",x"c2",x"1e"),
  1600 => (x"c2",x"78",x"c0",x"48"),
  1601 => (x"c0",x"48",x"dc",x"e9"),
  1602 => (x"87",x"fc",x"fd",x"78"),
  1603 => (x"48",x"c0",x"87",x"e1"),
  1604 => (x"00",x"00",x"4f",x"26"),
  1605 => (x"00",x"00",x"00",x"01"),
  1606 => (x"78",x"45",x"20",x"80"),
  1607 => (x"80",x"00",x"74",x"69"),
  1608 => (x"63",x"61",x"42",x"20"),
  1609 => (x"10",x"37",x"00",x"6b"),
  1610 => (x"2a",x"88",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"10",x"37",x"00"),
  1613 => (x"00",x"2a",x"a6",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"10",x"37"),
  1616 => (x"00",x"00",x"2a",x"c4"),
  1617 => (x"37",x"00",x"00",x"00"),
  1618 => (x"e2",x"00",x"00",x"10"),
  1619 => (x"00",x"00",x"00",x"2a"),
  1620 => (x"10",x"37",x"00",x"00"),
  1621 => (x"2b",x"00",x"00",x"00"),
  1622 => (x"00",x"00",x"00",x"00"),
  1623 => (x"00",x"10",x"37",x"00"),
  1624 => (x"00",x"2b",x"1e",x"00"),
  1625 => (x"00",x"00",x"00",x"00"),
  1626 => (x"00",x"00",x"10",x"37"),
  1627 => (x"00",x"00",x"2b",x"3c"),
  1628 => (x"74",x"00",x"00",x"00"),
  1629 => (x"00",x"00",x"00",x"12"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"13",x"44",x"00",x"00"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"f0",x"fe",x"1e",x"00"),
  1635 => (x"cd",x"78",x"c0",x"48"),
  1636 => (x"26",x"09",x"79",x"09"),
  1637 => (x"fe",x"1e",x"1e",x"4f"),
  1638 => (x"48",x"7e",x"bf",x"f0"),
  1639 => (x"1e",x"4f",x"26",x"26"),
  1640 => (x"c1",x"48",x"f0",x"fe"),
  1641 => (x"1e",x"4f",x"26",x"78"),
  1642 => (x"c0",x"48",x"f0",x"fe"),
  1643 => (x"1e",x"4f",x"26",x"78"),
  1644 => (x"52",x"c0",x"4a",x"71"),
  1645 => (x"0e",x"4f",x"26",x"52"),
  1646 => (x"5d",x"5c",x"5b",x"5e"),
  1647 => (x"71",x"86",x"f4",x"0e"),
  1648 => (x"7e",x"6d",x"97",x"4d"),
  1649 => (x"97",x"4c",x"a5",x"c1"),
  1650 => (x"a6",x"c8",x"48",x"6c"),
  1651 => (x"c4",x"48",x"6e",x"58"),
  1652 => (x"c5",x"05",x"a8",x"66"),
  1653 => (x"c0",x"48",x"ff",x"87"),
  1654 => (x"ca",x"ff",x"87",x"e6"),
  1655 => (x"49",x"a5",x"c2",x"87"),
  1656 => (x"71",x"4b",x"6c",x"97"),
  1657 => (x"6b",x"97",x"4b",x"a3"),
  1658 => (x"7e",x"6c",x"97",x"4b"),
  1659 => (x"80",x"c1",x"48",x"6e"),
  1660 => (x"c7",x"58",x"a6",x"c8"),
  1661 => (x"58",x"a6",x"cc",x"98"),
  1662 => (x"fe",x"7c",x"97",x"70"),
  1663 => (x"48",x"73",x"87",x"e1"),
  1664 => (x"4d",x"26",x"8e",x"f4"),
  1665 => (x"4b",x"26",x"4c",x"26"),
  1666 => (x"5e",x"0e",x"4f",x"26"),
  1667 => (x"f4",x"0e",x"5c",x"5b"),
  1668 => (x"d8",x"4c",x"71",x"86"),
  1669 => (x"ff",x"c3",x"4a",x"66"),
  1670 => (x"4b",x"a4",x"c2",x"9a"),
  1671 => (x"73",x"49",x"6c",x"97"),
  1672 => (x"51",x"72",x"49",x"a1"),
  1673 => (x"6e",x"7e",x"6c",x"97"),
  1674 => (x"c8",x"80",x"c1",x"48"),
  1675 => (x"98",x"c7",x"58",x"a6"),
  1676 => (x"70",x"58",x"a6",x"cc"),
  1677 => (x"ff",x"8e",x"f4",x"54"),
  1678 => (x"1e",x"1e",x"87",x"ca"),
  1679 => (x"e0",x"87",x"e8",x"fd"),
  1680 => (x"c0",x"49",x"4a",x"bf"),
  1681 => (x"02",x"99",x"c0",x"e0"),
  1682 => (x"1e",x"72",x"87",x"cb"),
  1683 => (x"49",x"da",x"ed",x"c2"),
  1684 => (x"c4",x"87",x"f7",x"fe"),
  1685 => (x"87",x"fd",x"fc",x"86"),
  1686 => (x"c2",x"fd",x"7e",x"70"),
  1687 => (x"4f",x"26",x"26",x"87"),
  1688 => (x"da",x"ed",x"c2",x"1e"),
  1689 => (x"87",x"c7",x"fd",x"49"),
  1690 => (x"49",x"fa",x"e8",x"c1"),
  1691 => (x"c2",x"87",x"da",x"fc"),
  1692 => (x"4f",x"26",x"87",x"fe"),
  1693 => (x"c2",x"1e",x"73",x"1e"),
  1694 => (x"fc",x"49",x"da",x"ed"),
  1695 => (x"4a",x"70",x"87",x"f9"),
  1696 => (x"04",x"aa",x"b7",x"c0"),
  1697 => (x"c3",x"87",x"cc",x"c2"),
  1698 => (x"c9",x"05",x"aa",x"f0"),
  1699 => (x"df",x"ec",x"c1",x"87"),
  1700 => (x"c1",x"78",x"c1",x"48"),
  1701 => (x"e0",x"c3",x"87",x"ed"),
  1702 => (x"87",x"c9",x"05",x"aa"),
  1703 => (x"48",x"e3",x"ec",x"c1"),
  1704 => (x"de",x"c1",x"78",x"c1"),
  1705 => (x"e3",x"ec",x"c1",x"87"),
  1706 => (x"87",x"c6",x"02",x"bf"),
  1707 => (x"4b",x"a2",x"c0",x"c2"),
  1708 => (x"4b",x"72",x"87",x"c2"),
  1709 => (x"bf",x"df",x"ec",x"c1"),
  1710 => (x"87",x"e0",x"c0",x"02"),
  1711 => (x"b7",x"c4",x"49",x"73"),
  1712 => (x"ed",x"c1",x"91",x"29"),
  1713 => (x"4a",x"73",x"81",x"ff"),
  1714 => (x"92",x"c2",x"9a",x"cf"),
  1715 => (x"30",x"72",x"48",x"c1"),
  1716 => (x"ba",x"ff",x"4a",x"70"),
  1717 => (x"98",x"69",x"48",x"72"),
  1718 => (x"87",x"db",x"79",x"70"),
  1719 => (x"b7",x"c4",x"49",x"73"),
  1720 => (x"ed",x"c1",x"91",x"29"),
  1721 => (x"4a",x"73",x"81",x"ff"),
  1722 => (x"92",x"c2",x"9a",x"cf"),
  1723 => (x"30",x"72",x"48",x"c3"),
  1724 => (x"69",x"48",x"4a",x"70"),
  1725 => (x"c1",x"79",x"70",x"b0"),
  1726 => (x"c0",x"48",x"e3",x"ec"),
  1727 => (x"df",x"ec",x"c1",x"78"),
  1728 => (x"c2",x"78",x"c0",x"48"),
  1729 => (x"fa",x"49",x"da",x"ed"),
  1730 => (x"4a",x"70",x"87",x"ed"),
  1731 => (x"03",x"aa",x"b7",x"c0"),
  1732 => (x"c0",x"87",x"f4",x"fd"),
  1733 => (x"26",x"87",x"c4",x"48"),
  1734 => (x"26",x"4c",x"26",x"4d"),
  1735 => (x"00",x"4f",x"26",x"4b"),
  1736 => (x"00",x"00",x"00",x"00"),
  1737 => (x"1e",x"00",x"00",x"00"),
  1738 => (x"fd",x"49",x"4a",x"71"),
  1739 => (x"4f",x"26",x"87",x"c6"),
  1740 => (x"72",x"4a",x"c0",x"1e"),
  1741 => (x"c1",x"91",x"c4",x"49"),
  1742 => (x"c0",x"81",x"ff",x"ed"),
  1743 => (x"d0",x"82",x"c1",x"79"),
  1744 => (x"ee",x"04",x"aa",x"b7"),
  1745 => (x"0e",x"4f",x"26",x"87"),
  1746 => (x"5d",x"5c",x"5b",x"5e"),
  1747 => (x"f9",x"4d",x"71",x"0e"),
  1748 => (x"4a",x"75",x"87",x"d5"),
  1749 => (x"92",x"2a",x"b7",x"c4"),
  1750 => (x"82",x"ff",x"ed",x"c1"),
  1751 => (x"9c",x"cf",x"4c",x"75"),
  1752 => (x"49",x"6a",x"94",x"c2"),
  1753 => (x"c3",x"2b",x"74",x"4b"),
  1754 => (x"74",x"48",x"c2",x"9b"),
  1755 => (x"ff",x"4c",x"70",x"30"),
  1756 => (x"71",x"48",x"74",x"bc"),
  1757 => (x"f8",x"7a",x"70",x"98"),
  1758 => (x"48",x"73",x"87",x"e5"),
  1759 => (x"00",x"87",x"d8",x"fe"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"1e",x"00",x"00",x"00"),
  1776 => (x"c8",x"48",x"d0",x"ff"),
  1777 => (x"48",x"71",x"78",x"e1"),
  1778 => (x"78",x"08",x"d4",x"ff"),
  1779 => (x"ff",x"1e",x"4f",x"26"),
  1780 => (x"e1",x"c8",x"48",x"d0"),
  1781 => (x"ff",x"48",x"71",x"78"),
  1782 => (x"c4",x"78",x"08",x"d4"),
  1783 => (x"d4",x"ff",x"48",x"66"),
  1784 => (x"4f",x"26",x"78",x"08"),
  1785 => (x"c4",x"4a",x"71",x"1e"),
  1786 => (x"72",x"1e",x"49",x"66"),
  1787 => (x"87",x"de",x"ff",x"49"),
  1788 => (x"c0",x"48",x"d0",x"ff"),
  1789 => (x"26",x"26",x"78",x"e0"),
  1790 => (x"1e",x"73",x"1e",x"4f"),
  1791 => (x"66",x"c8",x"4b",x"71"),
  1792 => (x"4a",x"73",x"1e",x"49"),
  1793 => (x"49",x"a2",x"e0",x"c1"),
  1794 => (x"26",x"87",x"d9",x"ff"),
  1795 => (x"4d",x"26",x"87",x"c4"),
  1796 => (x"4b",x"26",x"4c",x"26"),
  1797 => (x"ff",x"1e",x"4f",x"26"),
  1798 => (x"ff",x"c3",x"4a",x"d4"),
  1799 => (x"48",x"d0",x"ff",x"7a"),
  1800 => (x"de",x"78",x"e1",x"c0"),
  1801 => (x"e4",x"ed",x"c2",x"7a"),
  1802 => (x"48",x"49",x"7a",x"bf"),
  1803 => (x"7a",x"70",x"28",x"c8"),
  1804 => (x"28",x"d0",x"48",x"71"),
  1805 => (x"48",x"71",x"7a",x"70"),
  1806 => (x"7a",x"70",x"28",x"d8"),
  1807 => (x"c0",x"48",x"d0",x"ff"),
  1808 => (x"4f",x"26",x"78",x"e0"),
  1809 => (x"48",x"d0",x"ff",x"1e"),
  1810 => (x"71",x"78",x"c9",x"c8"),
  1811 => (x"08",x"d4",x"ff",x"48"),
  1812 => (x"1e",x"4f",x"26",x"78"),
  1813 => (x"eb",x"49",x"4a",x"71"),
  1814 => (x"48",x"d0",x"ff",x"87"),
  1815 => (x"4f",x"26",x"78",x"c8"),
  1816 => (x"71",x"1e",x"73",x"1e"),
  1817 => (x"f4",x"ed",x"c2",x"4b"),
  1818 => (x"87",x"c3",x"02",x"bf"),
  1819 => (x"ff",x"87",x"eb",x"c2"),
  1820 => (x"c9",x"c8",x"48",x"d0"),
  1821 => (x"c0",x"49",x"73",x"78"),
  1822 => (x"d4",x"ff",x"b1",x"e0"),
  1823 => (x"c2",x"78",x"71",x"48"),
  1824 => (x"c0",x"48",x"e8",x"ed"),
  1825 => (x"02",x"66",x"c8",x"78"),
  1826 => (x"ff",x"c3",x"87",x"c5"),
  1827 => (x"c0",x"87",x"c2",x"49"),
  1828 => (x"f0",x"ed",x"c2",x"49"),
  1829 => (x"02",x"66",x"cc",x"59"),
  1830 => (x"d5",x"c5",x"87",x"c6"),
  1831 => (x"87",x"c4",x"4a",x"d5"),
  1832 => (x"4a",x"ff",x"ff",x"cf"),
  1833 => (x"5a",x"f4",x"ed",x"c2"),
  1834 => (x"48",x"f4",x"ed",x"c2"),
  1835 => (x"87",x"c4",x"78",x"c1"),
  1836 => (x"4c",x"26",x"4d",x"26"),
  1837 => (x"4f",x"26",x"4b",x"26"),
  1838 => (x"5c",x"5b",x"5e",x"0e"),
  1839 => (x"4a",x"71",x"0e",x"5d"),
  1840 => (x"bf",x"f0",x"ed",x"c2"),
  1841 => (x"02",x"9a",x"72",x"4c"),
  1842 => (x"c8",x"49",x"87",x"cb"),
  1843 => (x"d6",x"f1",x"c1",x"91"),
  1844 => (x"c4",x"83",x"71",x"4b"),
  1845 => (x"d6",x"f5",x"c1",x"87"),
  1846 => (x"13",x"4d",x"c0",x"4b"),
  1847 => (x"c2",x"99",x"74",x"49"),
  1848 => (x"b9",x"bf",x"ec",x"ed"),
  1849 => (x"71",x"48",x"d4",x"ff"),
  1850 => (x"2c",x"b7",x"c1",x"78"),
  1851 => (x"ad",x"b7",x"c8",x"85"),
  1852 => (x"c2",x"87",x"e8",x"04"),
  1853 => (x"48",x"bf",x"e8",x"ed"),
  1854 => (x"ed",x"c2",x"80",x"c8"),
  1855 => (x"ef",x"fe",x"58",x"ec"),
  1856 => (x"1e",x"73",x"1e",x"87"),
  1857 => (x"4a",x"13",x"4b",x"71"),
  1858 => (x"87",x"cb",x"02",x"9a"),
  1859 => (x"e7",x"fe",x"49",x"72"),
  1860 => (x"9a",x"4a",x"13",x"87"),
  1861 => (x"fe",x"87",x"f5",x"05"),
  1862 => (x"c2",x"1e",x"87",x"da"),
  1863 => (x"49",x"bf",x"e8",x"ed"),
  1864 => (x"48",x"e8",x"ed",x"c2"),
  1865 => (x"c4",x"78",x"a1",x"c1"),
  1866 => (x"03",x"a9",x"b7",x"c0"),
  1867 => (x"d4",x"ff",x"87",x"db"),
  1868 => (x"ec",x"ed",x"c2",x"48"),
  1869 => (x"ed",x"c2",x"78",x"bf"),
  1870 => (x"c2",x"49",x"bf",x"e8"),
  1871 => (x"c1",x"48",x"e8",x"ed"),
  1872 => (x"c0",x"c4",x"78",x"a1"),
  1873 => (x"e5",x"04",x"a9",x"b7"),
  1874 => (x"48",x"d0",x"ff",x"87"),
  1875 => (x"ed",x"c2",x"78",x"c8"),
  1876 => (x"78",x"c0",x"48",x"f4"),
  1877 => (x"00",x"00",x"4f",x"26"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"5f",x"5f",x"00"),
  1881 => (x"03",x"00",x"00",x"00"),
  1882 => (x"03",x"03",x"00",x"03"),
  1883 => (x"7f",x"14",x"00",x"00"),
  1884 => (x"7f",x"7f",x"14",x"7f"),
  1885 => (x"24",x"00",x"00",x"14"),
  1886 => (x"3a",x"6b",x"6b",x"2e"),
  1887 => (x"6a",x"4c",x"00",x"12"),
  1888 => (x"56",x"6c",x"18",x"36"),
  1889 => (x"7e",x"30",x"00",x"32"),
  1890 => (x"3a",x"77",x"59",x"4f"),
  1891 => (x"00",x"00",x"40",x"68"),
  1892 => (x"00",x"03",x"07",x"04"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"41",x"63",x"3e",x"1c"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"1c",x"3e",x"63",x"41"),
  1897 => (x"2a",x"08",x"00",x"00"),
  1898 => (x"3e",x"1c",x"1c",x"3e"),
  1899 => (x"08",x"00",x"08",x"2a"),
  1900 => (x"08",x"3e",x"3e",x"08"),
  1901 => (x"00",x"00",x"00",x"08"),
  1902 => (x"00",x"60",x"e0",x"80"),
  1903 => (x"08",x"00",x"00",x"00"),
  1904 => (x"08",x"08",x"08",x"08"),
  1905 => (x"00",x"00",x"00",x"08"),
  1906 => (x"00",x"60",x"60",x"00"),
  1907 => (x"60",x"40",x"00",x"00"),
  1908 => (x"06",x"0c",x"18",x"30"),
  1909 => (x"3e",x"00",x"01",x"03"),
  1910 => (x"7f",x"4d",x"59",x"7f"),
  1911 => (x"04",x"00",x"00",x"3e"),
  1912 => (x"00",x"7f",x"7f",x"06"),
  1913 => (x"42",x"00",x"00",x"00"),
  1914 => (x"4f",x"59",x"71",x"63"),
  1915 => (x"22",x"00",x"00",x"46"),
  1916 => (x"7f",x"49",x"49",x"63"),
  1917 => (x"1c",x"18",x"00",x"36"),
  1918 => (x"7f",x"7f",x"13",x"16"),
  1919 => (x"27",x"00",x"00",x"10"),
  1920 => (x"7d",x"45",x"45",x"67"),
  1921 => (x"3c",x"00",x"00",x"39"),
  1922 => (x"79",x"49",x"4b",x"7e"),
  1923 => (x"01",x"00",x"00",x"30"),
  1924 => (x"0f",x"79",x"71",x"01"),
  1925 => (x"36",x"00",x"00",x"07"),
  1926 => (x"7f",x"49",x"49",x"7f"),
  1927 => (x"06",x"00",x"00",x"36"),
  1928 => (x"3f",x"69",x"49",x"4f"),
  1929 => (x"00",x"00",x"00",x"1e"),
  1930 => (x"00",x"66",x"66",x"00"),
  1931 => (x"00",x"00",x"00",x"00"),
  1932 => (x"00",x"66",x"e6",x"80"),
  1933 => (x"08",x"00",x"00",x"00"),
  1934 => (x"22",x"14",x"14",x"08"),
  1935 => (x"14",x"00",x"00",x"22"),
  1936 => (x"14",x"14",x"14",x"14"),
  1937 => (x"22",x"00",x"00",x"14"),
  1938 => (x"08",x"14",x"14",x"22"),
  1939 => (x"02",x"00",x"00",x"08"),
  1940 => (x"0f",x"59",x"51",x"03"),
  1941 => (x"7f",x"3e",x"00",x"06"),
  1942 => (x"1f",x"55",x"5d",x"41"),
  1943 => (x"7e",x"00",x"00",x"1e"),
  1944 => (x"7f",x"09",x"09",x"7f"),
  1945 => (x"7f",x"00",x"00",x"7e"),
  1946 => (x"7f",x"49",x"49",x"7f"),
  1947 => (x"1c",x"00",x"00",x"36"),
  1948 => (x"41",x"41",x"63",x"3e"),
  1949 => (x"7f",x"00",x"00",x"41"),
  1950 => (x"3e",x"63",x"41",x"7f"),
  1951 => (x"7f",x"00",x"00",x"1c"),
  1952 => (x"41",x"49",x"49",x"7f"),
  1953 => (x"7f",x"00",x"00",x"41"),
  1954 => (x"01",x"09",x"09",x"7f"),
  1955 => (x"3e",x"00",x"00",x"01"),
  1956 => (x"7b",x"49",x"41",x"7f"),
  1957 => (x"7f",x"00",x"00",x"7a"),
  1958 => (x"7f",x"08",x"08",x"7f"),
  1959 => (x"00",x"00",x"00",x"7f"),
  1960 => (x"41",x"7f",x"7f",x"41"),
  1961 => (x"20",x"00",x"00",x"00"),
  1962 => (x"7f",x"40",x"40",x"60"),
  1963 => (x"7f",x"7f",x"00",x"3f"),
  1964 => (x"63",x"36",x"1c",x"08"),
  1965 => (x"7f",x"00",x"00",x"41"),
  1966 => (x"40",x"40",x"40",x"7f"),
  1967 => (x"7f",x"7f",x"00",x"40"),
  1968 => (x"7f",x"06",x"0c",x"06"),
  1969 => (x"7f",x"7f",x"00",x"7f"),
  1970 => (x"7f",x"18",x"0c",x"06"),
  1971 => (x"3e",x"00",x"00",x"7f"),
  1972 => (x"7f",x"41",x"41",x"7f"),
  1973 => (x"7f",x"00",x"00",x"3e"),
  1974 => (x"0f",x"09",x"09",x"7f"),
  1975 => (x"7f",x"3e",x"00",x"06"),
  1976 => (x"7e",x"7f",x"61",x"41"),
  1977 => (x"7f",x"00",x"00",x"40"),
  1978 => (x"7f",x"19",x"09",x"7f"),
  1979 => (x"26",x"00",x"00",x"66"),
  1980 => (x"7b",x"59",x"4d",x"6f"),
  1981 => (x"01",x"00",x"00",x"32"),
  1982 => (x"01",x"7f",x"7f",x"01"),
  1983 => (x"3f",x"00",x"00",x"01"),
  1984 => (x"7f",x"40",x"40",x"7f"),
  1985 => (x"0f",x"00",x"00",x"3f"),
  1986 => (x"3f",x"70",x"70",x"3f"),
  1987 => (x"7f",x"7f",x"00",x"0f"),
  1988 => (x"7f",x"30",x"18",x"30"),
  1989 => (x"63",x"41",x"00",x"7f"),
  1990 => (x"36",x"1c",x"1c",x"36"),
  1991 => (x"03",x"01",x"41",x"63"),
  1992 => (x"06",x"7c",x"7c",x"06"),
  1993 => (x"71",x"61",x"01",x"03"),
  1994 => (x"43",x"47",x"4d",x"59"),
  1995 => (x"00",x"00",x"00",x"41"),
  1996 => (x"41",x"41",x"7f",x"7f"),
  1997 => (x"03",x"01",x"00",x"00"),
  1998 => (x"30",x"18",x"0c",x"06"),
  1999 => (x"00",x"00",x"40",x"60"),
  2000 => (x"7f",x"7f",x"41",x"41"),
  2001 => (x"0c",x"08",x"00",x"00"),
  2002 => (x"0c",x"06",x"03",x"06"),
  2003 => (x"80",x"80",x"00",x"08"),
  2004 => (x"80",x"80",x"80",x"80"),
  2005 => (x"00",x"00",x"00",x"80"),
  2006 => (x"04",x"07",x"03",x"00"),
  2007 => (x"20",x"00",x"00",x"00"),
  2008 => (x"7c",x"54",x"54",x"74"),
  2009 => (x"7f",x"00",x"00",x"78"),
  2010 => (x"7c",x"44",x"44",x"7f"),
  2011 => (x"38",x"00",x"00",x"38"),
  2012 => (x"44",x"44",x"44",x"7c"),
  2013 => (x"38",x"00",x"00",x"00"),
  2014 => (x"7f",x"44",x"44",x"7c"),
  2015 => (x"38",x"00",x"00",x"7f"),
  2016 => (x"5c",x"54",x"54",x"7c"),
  2017 => (x"04",x"00",x"00",x"18"),
  2018 => (x"05",x"05",x"7f",x"7e"),
  2019 => (x"18",x"00",x"00",x"00"),
  2020 => (x"fc",x"a4",x"a4",x"bc"),
  2021 => (x"7f",x"00",x"00",x"7c"),
  2022 => (x"7c",x"04",x"04",x"7f"),
  2023 => (x"00",x"00",x"00",x"78"),
  2024 => (x"40",x"7d",x"3d",x"00"),
  2025 => (x"80",x"00",x"00",x"00"),
  2026 => (x"7d",x"fd",x"80",x"80"),
  2027 => (x"7f",x"00",x"00",x"00"),
  2028 => (x"6c",x"38",x"10",x"7f"),
  2029 => (x"00",x"00",x"00",x"44"),
  2030 => (x"40",x"7f",x"3f",x"00"),
  2031 => (x"7c",x"7c",x"00",x"00"),
  2032 => (x"7c",x"0c",x"18",x"0c"),
  2033 => (x"7c",x"00",x"00",x"78"),
  2034 => (x"7c",x"04",x"04",x"7c"),
  2035 => (x"38",x"00",x"00",x"78"),
  2036 => (x"7c",x"44",x"44",x"7c"),
  2037 => (x"fc",x"00",x"00",x"38"),
  2038 => (x"3c",x"24",x"24",x"fc"),
  2039 => (x"18",x"00",x"00",x"18"),
  2040 => (x"fc",x"24",x"24",x"3c"),
  2041 => (x"7c",x"00",x"00",x"fc"),
  2042 => (x"0c",x"04",x"04",x"7c"),
  2043 => (x"48",x"00",x"00",x"08"),
  2044 => (x"74",x"54",x"54",x"5c"),
  2045 => (x"04",x"00",x"00",x"20"),
  2046 => (x"44",x"44",x"7f",x"3f"),
  2047 => (x"3c",x"00",x"00",x"00"),
  2048 => (x"7c",x"40",x"40",x"7c"),
  2049 => (x"1c",x"00",x"00",x"7c"),
  2050 => (x"3c",x"60",x"60",x"3c"),
  2051 => (x"7c",x"3c",x"00",x"1c"),
  2052 => (x"7c",x"60",x"30",x"60"),
  2053 => (x"6c",x"44",x"00",x"3c"),
  2054 => (x"6c",x"38",x"10",x"38"),
  2055 => (x"1c",x"00",x"00",x"44"),
  2056 => (x"3c",x"60",x"e0",x"bc"),
  2057 => (x"44",x"00",x"00",x"1c"),
  2058 => (x"4c",x"5c",x"74",x"64"),
  2059 => (x"08",x"00",x"00",x"44"),
  2060 => (x"41",x"77",x"3e",x"08"),
  2061 => (x"00",x"00",x"00",x"41"),
  2062 => (x"00",x"7f",x"7f",x"00"),
  2063 => (x"41",x"00",x"00",x"00"),
  2064 => (x"08",x"3e",x"77",x"41"),
  2065 => (x"01",x"02",x"00",x"08"),
  2066 => (x"02",x"02",x"03",x"01"),
  2067 => (x"7f",x"7f",x"00",x"01"),
  2068 => (x"7f",x"7f",x"7f",x"7f"),
  2069 => (x"08",x"08",x"00",x"7f"),
  2070 => (x"3e",x"3e",x"1c",x"1c"),
  2071 => (x"7f",x"7f",x"7f",x"7f"),
  2072 => (x"1c",x"1c",x"3e",x"3e"),
  2073 => (x"10",x"00",x"08",x"08"),
  2074 => (x"18",x"7c",x"7c",x"18"),
  2075 => (x"10",x"00",x"00",x"10"),
  2076 => (x"30",x"7c",x"7c",x"30"),
  2077 => (x"30",x"10",x"00",x"10"),
  2078 => (x"1e",x"78",x"60",x"60"),
  2079 => (x"66",x"42",x"00",x"06"),
  2080 => (x"66",x"3c",x"18",x"3c"),
  2081 => (x"38",x"78",x"00",x"42"),
  2082 => (x"6c",x"c6",x"c2",x"6a"),
  2083 => (x"00",x"60",x"00",x"38"),
  2084 => (x"00",x"00",x"60",x"00"),
  2085 => (x"5e",x"0e",x"00",x"60"),
  2086 => (x"0e",x"5d",x"5c",x"5b"),
  2087 => (x"c2",x"4c",x"71",x"1e"),
  2088 => (x"4d",x"bf",x"c5",x"ee"),
  2089 => (x"1e",x"c0",x"4b",x"c0"),
  2090 => (x"c7",x"02",x"ab",x"74"),
  2091 => (x"48",x"a6",x"c4",x"87"),
  2092 => (x"87",x"c5",x"78",x"c0"),
  2093 => (x"c1",x"48",x"a6",x"c4"),
  2094 => (x"1e",x"66",x"c4",x"78"),
  2095 => (x"df",x"ee",x"49",x"73"),
  2096 => (x"c0",x"86",x"c8",x"87"),
  2097 => (x"ef",x"ef",x"49",x"e0"),
  2098 => (x"4a",x"a5",x"c4",x"87"),
  2099 => (x"f0",x"f0",x"49",x"6a"),
  2100 => (x"87",x"c6",x"f1",x"87"),
  2101 => (x"83",x"c1",x"85",x"cb"),
  2102 => (x"04",x"ab",x"b7",x"c8"),
  2103 => (x"26",x"87",x"c7",x"ff"),
  2104 => (x"4c",x"26",x"4d",x"26"),
  2105 => (x"4f",x"26",x"4b",x"26"),
  2106 => (x"c2",x"4a",x"71",x"1e"),
  2107 => (x"c2",x"5a",x"c9",x"ee"),
  2108 => (x"c7",x"48",x"c9",x"ee"),
  2109 => (x"dd",x"fe",x"49",x"78"),
  2110 => (x"1e",x"4f",x"26",x"87"),
  2111 => (x"4a",x"71",x"1e",x"73"),
  2112 => (x"03",x"aa",x"b7",x"c0"),
  2113 => (x"d2",x"c2",x"87",x"d3"),
  2114 => (x"c4",x"05",x"bf",x"ee"),
  2115 => (x"c2",x"4b",x"c1",x"87"),
  2116 => (x"c2",x"4b",x"c0",x"87"),
  2117 => (x"c4",x"5b",x"f2",x"d2"),
  2118 => (x"f2",x"d2",x"c2",x"87"),
  2119 => (x"ee",x"d2",x"c2",x"5a"),
  2120 => (x"9a",x"c1",x"4a",x"bf"),
  2121 => (x"49",x"a2",x"c0",x"c1"),
  2122 => (x"fc",x"87",x"e8",x"ec"),
  2123 => (x"ee",x"d2",x"c2",x"48"),
  2124 => (x"ef",x"fe",x"78",x"bf"),
  2125 => (x"4a",x"71",x"1e",x"87"),
  2126 => (x"72",x"1e",x"66",x"c4"),
  2127 => (x"87",x"f9",x"ea",x"49"),
  2128 => (x"1e",x"4f",x"26",x"26"),
  2129 => (x"d4",x"ff",x"4a",x"71"),
  2130 => (x"78",x"ff",x"c3",x"48"),
  2131 => (x"c0",x"48",x"d0",x"ff"),
  2132 => (x"d4",x"ff",x"78",x"e1"),
  2133 => (x"72",x"78",x"c1",x"48"),
  2134 => (x"71",x"31",x"c4",x"49"),
  2135 => (x"48",x"d0",x"ff",x"78"),
  2136 => (x"26",x"78",x"e0",x"c0"),
  2137 => (x"d2",x"c2",x"1e",x"4f"),
  2138 => (x"e6",x"49",x"bf",x"ee"),
  2139 => (x"ed",x"c2",x"87",x"f9"),
  2140 => (x"bf",x"e8",x"48",x"fd"),
  2141 => (x"f9",x"ed",x"c2",x"78"),
  2142 => (x"78",x"bf",x"ec",x"48"),
  2143 => (x"bf",x"fd",x"ed",x"c2"),
  2144 => (x"ff",x"c3",x"49",x"4a"),
  2145 => (x"2a",x"b7",x"c8",x"99"),
  2146 => (x"b0",x"71",x"48",x"72"),
  2147 => (x"58",x"c5",x"ee",x"c2"),
  2148 => (x"5e",x"0e",x"4f",x"26"),
  2149 => (x"0e",x"5d",x"5c",x"5b"),
  2150 => (x"c8",x"ff",x"4b",x"71"),
  2151 => (x"f8",x"ed",x"c2",x"87"),
  2152 => (x"73",x"50",x"c0",x"48"),
  2153 => (x"87",x"df",x"e6",x"49"),
  2154 => (x"c2",x"4c",x"49",x"70"),
  2155 => (x"49",x"ee",x"cb",x"9c"),
  2156 => (x"70",x"87",x"c3",x"cc"),
  2157 => (x"ed",x"c2",x"4d",x"49"),
  2158 => (x"05",x"bf",x"97",x"f8"),
  2159 => (x"d0",x"87",x"e2",x"c1"),
  2160 => (x"ee",x"c2",x"49",x"66"),
  2161 => (x"05",x"99",x"bf",x"c1"),
  2162 => (x"66",x"d4",x"87",x"d6"),
  2163 => (x"f9",x"ed",x"c2",x"49"),
  2164 => (x"cb",x"05",x"99",x"bf"),
  2165 => (x"e5",x"49",x"73",x"87"),
  2166 => (x"98",x"70",x"87",x"ed"),
  2167 => (x"87",x"c1",x"c1",x"02"),
  2168 => (x"c0",x"fe",x"4c",x"c1"),
  2169 => (x"cb",x"49",x"75",x"87"),
  2170 => (x"98",x"70",x"87",x"d8"),
  2171 => (x"c2",x"87",x"c6",x"02"),
  2172 => (x"c1",x"48",x"f8",x"ed"),
  2173 => (x"f8",x"ed",x"c2",x"50"),
  2174 => (x"c0",x"05",x"bf",x"97"),
  2175 => (x"ee",x"c2",x"87",x"e3"),
  2176 => (x"d0",x"49",x"bf",x"c1"),
  2177 => (x"ff",x"05",x"99",x"66"),
  2178 => (x"ed",x"c2",x"87",x"d6"),
  2179 => (x"d4",x"49",x"bf",x"f9"),
  2180 => (x"ff",x"05",x"99",x"66"),
  2181 => (x"49",x"73",x"87",x"ca"),
  2182 => (x"70",x"87",x"ec",x"e4"),
  2183 => (x"ff",x"fe",x"05",x"98"),
  2184 => (x"fa",x"48",x"74",x"87"),
  2185 => (x"5e",x"0e",x"87",x"fa"),
  2186 => (x"0e",x"5d",x"5c",x"5b"),
  2187 => (x"4d",x"c0",x"86",x"f8"),
  2188 => (x"7e",x"bf",x"ec",x"4c"),
  2189 => (x"c2",x"48",x"a6",x"c4"),
  2190 => (x"78",x"bf",x"c5",x"ee"),
  2191 => (x"1e",x"c0",x"1e",x"c1"),
  2192 => (x"cd",x"fd",x"49",x"c7"),
  2193 => (x"70",x"86",x"c8",x"87"),
  2194 => (x"87",x"cd",x"02",x"98"),
  2195 => (x"ea",x"fa",x"49",x"ff"),
  2196 => (x"49",x"da",x"c1",x"87"),
  2197 => (x"c1",x"87",x"f0",x"e3"),
  2198 => (x"f8",x"ed",x"c2",x"4d"),
  2199 => (x"cf",x"02",x"bf",x"97"),
  2200 => (x"e6",x"d2",x"c2",x"87"),
  2201 => (x"b9",x"c1",x"49",x"bf"),
  2202 => (x"59",x"ea",x"d2",x"c2"),
  2203 => (x"87",x"d3",x"fb",x"71"),
  2204 => (x"bf",x"fd",x"ed",x"c2"),
  2205 => (x"ee",x"d2",x"c2",x"4b"),
  2206 => (x"d9",x"c1",x"05",x"bf"),
  2207 => (x"48",x"a6",x"c4",x"87"),
  2208 => (x"78",x"c0",x"c0",x"c8"),
  2209 => (x"7e",x"e1",x"db",x"c2"),
  2210 => (x"49",x"bf",x"97",x"6e"),
  2211 => (x"80",x"c1",x"48",x"6e"),
  2212 => (x"e2",x"71",x"7e",x"70"),
  2213 => (x"98",x"70",x"87",x"f1"),
  2214 => (x"c4",x"87",x"c3",x"02"),
  2215 => (x"66",x"c4",x"b3",x"66"),
  2216 => (x"28",x"b7",x"c1",x"48"),
  2217 => (x"70",x"58",x"a6",x"c8"),
  2218 => (x"db",x"ff",x"05",x"98"),
  2219 => (x"49",x"fd",x"c3",x"87"),
  2220 => (x"c3",x"87",x"d4",x"e2"),
  2221 => (x"ce",x"e2",x"49",x"fa"),
  2222 => (x"c3",x"49",x"73",x"87"),
  2223 => (x"1e",x"71",x"99",x"ff"),
  2224 => (x"f0",x"f9",x"49",x"c0"),
  2225 => (x"c8",x"49",x"73",x"87"),
  2226 => (x"1e",x"71",x"29",x"b7"),
  2227 => (x"e4",x"f9",x"49",x"c1"),
  2228 => (x"c5",x"86",x"c8",x"87"),
  2229 => (x"ee",x"c2",x"87",x"fa"),
  2230 => (x"9b",x"4b",x"bf",x"c1"),
  2231 => (x"c2",x"87",x"dd",x"02"),
  2232 => (x"49",x"bf",x"ea",x"d2"),
  2233 => (x"70",x"87",x"db",x"c7"),
  2234 => (x"87",x"c4",x"05",x"98"),
  2235 => (x"87",x"d2",x"4b",x"c0"),
  2236 => (x"c7",x"49",x"e0",x"c2"),
  2237 => (x"d2",x"c2",x"87",x"c0"),
  2238 => (x"87",x"c6",x"58",x"ee"),
  2239 => (x"48",x"ea",x"d2",x"c2"),
  2240 => (x"49",x"73",x"78",x"c0"),
  2241 => (x"ce",x"05",x"99",x"c2"),
  2242 => (x"49",x"eb",x"c3",x"87"),
  2243 => (x"70",x"87",x"f8",x"e0"),
  2244 => (x"02",x"99",x"c2",x"49"),
  2245 => (x"fb",x"87",x"c2",x"c0"),
  2246 => (x"c1",x"49",x"73",x"4c"),
  2247 => (x"87",x"ce",x"05",x"99"),
  2248 => (x"e0",x"49",x"f4",x"c3"),
  2249 => (x"49",x"70",x"87",x"e1"),
  2250 => (x"c0",x"02",x"99",x"c2"),
  2251 => (x"4c",x"fa",x"87",x"c2"),
  2252 => (x"99",x"c8",x"49",x"73"),
  2253 => (x"c3",x"87",x"cd",x"05"),
  2254 => (x"ca",x"e0",x"49",x"f5"),
  2255 => (x"c2",x"49",x"70",x"87"),
  2256 => (x"87",x"d6",x"02",x"99"),
  2257 => (x"bf",x"c9",x"ee",x"c2"),
  2258 => (x"87",x"ca",x"c0",x"02"),
  2259 => (x"c2",x"88",x"c1",x"48"),
  2260 => (x"c0",x"58",x"cd",x"ee"),
  2261 => (x"4c",x"ff",x"87",x"c2"),
  2262 => (x"49",x"73",x"4d",x"c1"),
  2263 => (x"c0",x"05",x"99",x"c4"),
  2264 => (x"f2",x"c3",x"87",x"ce"),
  2265 => (x"de",x"df",x"ff",x"49"),
  2266 => (x"c2",x"49",x"70",x"87"),
  2267 => (x"87",x"dc",x"02",x"99"),
  2268 => (x"bf",x"c9",x"ee",x"c2"),
  2269 => (x"b7",x"c7",x"48",x"7e"),
  2270 => (x"cb",x"c0",x"03",x"a8"),
  2271 => (x"c1",x"48",x"6e",x"87"),
  2272 => (x"cd",x"ee",x"c2",x"80"),
  2273 => (x"87",x"c2",x"c0",x"58"),
  2274 => (x"4d",x"c1",x"4c",x"fe"),
  2275 => (x"ff",x"49",x"fd",x"c3"),
  2276 => (x"70",x"87",x"f4",x"de"),
  2277 => (x"02",x"99",x"c2",x"49"),
  2278 => (x"c2",x"87",x"d5",x"c0"),
  2279 => (x"02",x"bf",x"c9",x"ee"),
  2280 => (x"c2",x"87",x"c9",x"c0"),
  2281 => (x"c0",x"48",x"c9",x"ee"),
  2282 => (x"87",x"c2",x"c0",x"78"),
  2283 => (x"4d",x"c1",x"4c",x"fd"),
  2284 => (x"ff",x"49",x"fa",x"c3"),
  2285 => (x"70",x"87",x"d0",x"de"),
  2286 => (x"02",x"99",x"c2",x"49"),
  2287 => (x"c2",x"87",x"d9",x"c0"),
  2288 => (x"48",x"bf",x"c9",x"ee"),
  2289 => (x"03",x"a8",x"b7",x"c7"),
  2290 => (x"c2",x"87",x"c9",x"c0"),
  2291 => (x"c7",x"48",x"c9",x"ee"),
  2292 => (x"87",x"c2",x"c0",x"78"),
  2293 => (x"4d",x"c1",x"4c",x"fc"),
  2294 => (x"03",x"ac",x"b7",x"c0"),
  2295 => (x"c4",x"87",x"d3",x"c0"),
  2296 => (x"d8",x"c1",x"48",x"66"),
  2297 => (x"6e",x"7e",x"70",x"80"),
  2298 => (x"c5",x"c0",x"02",x"bf"),
  2299 => (x"49",x"74",x"4b",x"87"),
  2300 => (x"1e",x"c0",x"0f",x"73"),
  2301 => (x"c1",x"1e",x"f0",x"c3"),
  2302 => (x"d5",x"f6",x"49",x"da"),
  2303 => (x"70",x"86",x"c8",x"87"),
  2304 => (x"d8",x"c0",x"02",x"98"),
  2305 => (x"c9",x"ee",x"c2",x"87"),
  2306 => (x"49",x"6e",x"7e",x"bf"),
  2307 => (x"66",x"c4",x"91",x"cb"),
  2308 => (x"6a",x"82",x"71",x"4a"),
  2309 => (x"87",x"c5",x"c0",x"02"),
  2310 => (x"73",x"49",x"6e",x"4b"),
  2311 => (x"02",x"9d",x"75",x"0f"),
  2312 => (x"c2",x"87",x"c8",x"c0"),
  2313 => (x"49",x"bf",x"c9",x"ee"),
  2314 => (x"c2",x"87",x"eb",x"f1"),
  2315 => (x"02",x"bf",x"f2",x"d2"),
  2316 => (x"49",x"87",x"dd",x"c0"),
  2317 => (x"70",x"87",x"cb",x"c2"),
  2318 => (x"d3",x"c0",x"02",x"98"),
  2319 => (x"c9",x"ee",x"c2",x"87"),
  2320 => (x"d1",x"f1",x"49",x"bf"),
  2321 => (x"f2",x"49",x"c0",x"87"),
  2322 => (x"d2",x"c2",x"87",x"f1"),
  2323 => (x"78",x"c0",x"48",x"f2"),
  2324 => (x"cb",x"f2",x"8e",x"f8"),
  2325 => (x"5b",x"5e",x"0e",x"87"),
  2326 => (x"1e",x"0e",x"5d",x"5c"),
  2327 => (x"ee",x"c2",x"4c",x"71"),
  2328 => (x"c1",x"49",x"bf",x"c5"),
  2329 => (x"c1",x"4d",x"a1",x"cd"),
  2330 => (x"7e",x"69",x"81",x"d1"),
  2331 => (x"cf",x"02",x"9c",x"74"),
  2332 => (x"4b",x"a5",x"c4",x"87"),
  2333 => (x"ee",x"c2",x"7b",x"74"),
  2334 => (x"f1",x"49",x"bf",x"c5"),
  2335 => (x"7b",x"6e",x"87",x"ea"),
  2336 => (x"c4",x"05",x"9c",x"74"),
  2337 => (x"c2",x"4b",x"c0",x"87"),
  2338 => (x"73",x"4b",x"c1",x"87"),
  2339 => (x"87",x"eb",x"f1",x"49"),
  2340 => (x"c7",x"02",x"66",x"d4"),
  2341 => (x"87",x"de",x"49",x"87"),
  2342 => (x"87",x"c2",x"4a",x"70"),
  2343 => (x"d2",x"c2",x"4a",x"c0"),
  2344 => (x"f0",x"26",x"5a",x"f6"),
  2345 => (x"00",x"00",x"87",x"fa"),
  2346 => (x"00",x"00",x"00",x"00"),
  2347 => (x"00",x"00",x"00",x"00"),
  2348 => (x"00",x"00",x"00",x"00"),
  2349 => (x"71",x"1e",x"00",x"00"),
  2350 => (x"bf",x"c8",x"ff",x"4a"),
  2351 => (x"48",x"a1",x"72",x"49"),
  2352 => (x"ff",x"1e",x"4f",x"26"),
  2353 => (x"fe",x"89",x"bf",x"c8"),
  2354 => (x"c0",x"c0",x"c0",x"c0"),
  2355 => (x"c4",x"01",x"a9",x"c0"),
  2356 => (x"c2",x"4a",x"c0",x"87"),
  2357 => (x"72",x"4a",x"c1",x"87"),
  2358 => (x"0e",x"4f",x"26",x"48"),
  2359 => (x"5d",x"5c",x"5b",x"5e"),
  2360 => (x"ff",x"4b",x"71",x"0e"),
  2361 => (x"66",x"d0",x"4c",x"d4"),
  2362 => (x"d6",x"78",x"c0",x"48"),
  2363 => (x"ce",x"db",x"ff",x"49"),
  2364 => (x"7c",x"ff",x"c3",x"87"),
  2365 => (x"ff",x"c3",x"49",x"6c"),
  2366 => (x"49",x"4d",x"71",x"99"),
  2367 => (x"c1",x"99",x"f0",x"c3"),
  2368 => (x"cb",x"05",x"a9",x"e0"),
  2369 => (x"7c",x"ff",x"c3",x"87"),
  2370 => (x"98",x"c3",x"48",x"6c"),
  2371 => (x"78",x"08",x"66",x"d0"),
  2372 => (x"6c",x"7c",x"ff",x"c3"),
  2373 => (x"31",x"c8",x"49",x"4a"),
  2374 => (x"6c",x"7c",x"ff",x"c3"),
  2375 => (x"72",x"b2",x"71",x"4a"),
  2376 => (x"c3",x"31",x"c8",x"49"),
  2377 => (x"4a",x"6c",x"7c",x"ff"),
  2378 => (x"49",x"72",x"b2",x"71"),
  2379 => (x"ff",x"c3",x"31",x"c8"),
  2380 => (x"71",x"4a",x"6c",x"7c"),
  2381 => (x"48",x"d0",x"ff",x"b2"),
  2382 => (x"73",x"78",x"e0",x"c0"),
  2383 => (x"87",x"c2",x"02",x"9b"),
  2384 => (x"48",x"75",x"7b",x"72"),
  2385 => (x"4c",x"26",x"4d",x"26"),
  2386 => (x"4f",x"26",x"4b",x"26"),
  2387 => (x"0e",x"4f",x"26",x"1e"),
  2388 => (x"0e",x"5c",x"5b",x"5e"),
  2389 => (x"1e",x"76",x"86",x"f8"),
  2390 => (x"fd",x"49",x"a6",x"c8"),
  2391 => (x"86",x"c4",x"87",x"fd"),
  2392 => (x"48",x"6e",x"4b",x"70"),
  2393 => (x"c2",x"03",x"a8",x"c2"),
  2394 => (x"4a",x"73",x"87",x"f0"),
  2395 => (x"c1",x"9a",x"f0",x"c3"),
  2396 => (x"c7",x"02",x"aa",x"d0"),
  2397 => (x"aa",x"e0",x"c1",x"87"),
  2398 => (x"87",x"de",x"c2",x"05"),
  2399 => (x"99",x"c8",x"49",x"73"),
  2400 => (x"ff",x"87",x"c3",x"02"),
  2401 => (x"4c",x"73",x"87",x"c6"),
  2402 => (x"ac",x"c2",x"9c",x"c3"),
  2403 => (x"87",x"c2",x"c1",x"05"),
  2404 => (x"c9",x"49",x"66",x"c4"),
  2405 => (x"c4",x"1e",x"71",x"31"),
  2406 => (x"92",x"d4",x"4a",x"66"),
  2407 => (x"49",x"cd",x"ee",x"c2"),
  2408 => (x"d0",x"fe",x"81",x"72"),
  2409 => (x"49",x"d8",x"87",x"eb"),
  2410 => (x"87",x"d3",x"d8",x"ff"),
  2411 => (x"c2",x"1e",x"c0",x"c8"),
  2412 => (x"fd",x"49",x"ea",x"dc"),
  2413 => (x"ff",x"87",x"e7",x"ec"),
  2414 => (x"e0",x"c0",x"48",x"d0"),
  2415 => (x"ea",x"dc",x"c2",x"78"),
  2416 => (x"4a",x"66",x"cc",x"1e"),
  2417 => (x"ee",x"c2",x"92",x"d4"),
  2418 => (x"81",x"72",x"49",x"cd"),
  2419 => (x"87",x"f2",x"ce",x"fe"),
  2420 => (x"ac",x"c1",x"86",x"cc"),
  2421 => (x"87",x"c2",x"c1",x"05"),
  2422 => (x"c9",x"49",x"66",x"c4"),
  2423 => (x"c4",x"1e",x"71",x"31"),
  2424 => (x"92",x"d4",x"4a",x"66"),
  2425 => (x"49",x"cd",x"ee",x"c2"),
  2426 => (x"cf",x"fe",x"81",x"72"),
  2427 => (x"dc",x"c2",x"87",x"e3"),
  2428 => (x"66",x"c8",x"1e",x"ea"),
  2429 => (x"c2",x"92",x"d4",x"4a"),
  2430 => (x"72",x"49",x"cd",x"ee"),
  2431 => (x"f2",x"cc",x"fe",x"81"),
  2432 => (x"ff",x"49",x"d7",x"87"),
  2433 => (x"c8",x"87",x"f8",x"d6"),
  2434 => (x"dc",x"c2",x"1e",x"c0"),
  2435 => (x"ea",x"fd",x"49",x"ea"),
  2436 => (x"86",x"cc",x"87",x"e5"),
  2437 => (x"c0",x"48",x"d0",x"ff"),
  2438 => (x"8e",x"f8",x"78",x"e0"),
  2439 => (x"0e",x"87",x"e7",x"fc"),
  2440 => (x"5d",x"5c",x"5b",x"5e"),
  2441 => (x"4d",x"71",x"1e",x"0e"),
  2442 => (x"d4",x"4c",x"d4",x"ff"),
  2443 => (x"c3",x"48",x"7e",x"66"),
  2444 => (x"c5",x"06",x"a8",x"b7"),
  2445 => (x"c1",x"48",x"c0",x"87"),
  2446 => (x"49",x"75",x"87",x"e2"),
  2447 => (x"87",x"de",x"dd",x"fe"),
  2448 => (x"66",x"c4",x"1e",x"75"),
  2449 => (x"c2",x"93",x"d4",x"4b"),
  2450 => (x"73",x"83",x"cd",x"ee"),
  2451 => (x"ef",x"c6",x"fe",x"49"),
  2452 => (x"6b",x"83",x"c8",x"87"),
  2453 => (x"48",x"d0",x"ff",x"4b"),
  2454 => (x"dd",x"78",x"e1",x"c8"),
  2455 => (x"c3",x"49",x"73",x"7c"),
  2456 => (x"7c",x"71",x"99",x"ff"),
  2457 => (x"b7",x"c8",x"49",x"73"),
  2458 => (x"99",x"ff",x"c3",x"29"),
  2459 => (x"49",x"73",x"7c",x"71"),
  2460 => (x"c3",x"29",x"b7",x"d0"),
  2461 => (x"7c",x"71",x"99",x"ff"),
  2462 => (x"b7",x"d8",x"49",x"73"),
  2463 => (x"c0",x"7c",x"71",x"29"),
  2464 => (x"7c",x"7c",x"7c",x"7c"),
  2465 => (x"7c",x"7c",x"7c",x"7c"),
  2466 => (x"7c",x"7c",x"7c",x"7c"),
  2467 => (x"c4",x"78",x"e0",x"c0"),
  2468 => (x"49",x"dc",x"1e",x"66"),
  2469 => (x"87",x"cc",x"d5",x"ff"),
  2470 => (x"48",x"73",x"86",x"c8"),
  2471 => (x"87",x"e4",x"fa",x"26"),
  2472 => (x"c0",x"1e",x"73",x"1e"),
  2473 => (x"f5",x"db",x"c2",x"4b"),
  2474 => (x"c2",x"50",x"c0",x"48"),
  2475 => (x"49",x"bf",x"f1",x"db"),
  2476 => (x"87",x"ce",x"df",x"fe"),
  2477 => (x"c4",x"05",x"98",x"70"),
  2478 => (x"c9",x"db",x"c2",x"87"),
  2479 => (x"c4",x"48",x"73",x"4b"),
  2480 => (x"26",x"4d",x"26",x"87"),
  2481 => (x"26",x"4b",x"26",x"4c"),
  2482 => (x"6f",x"68",x"53",x"4f"),
  2483 => (x"69",x"68",x"2f",x"77"),
  2484 => (x"4f",x"20",x"65",x"64"),
  2485 => (x"3d",x"20",x"44",x"53"),
  2486 => (x"79",x"65",x"6b",x"20"),
  2487 => (x"32",x"31",x"46",x"20"),
  2488 => (x"14",x"12",x"58",x"00"),
  2489 => (x"1c",x"1b",x"1d",x"11"),
  2490 => (x"94",x"59",x"5a",x"23"),
  2491 => (x"eb",x"f2",x"f5",x"91"),
  2492 => (x"00",x"26",x"f6",x"f4"),
  2493 => (x"55",x"41",x"00",x"00"),
  2494 => (x"4f",x"42",x"4f",x"54"),
  2495 => (x"45",x"4e",x"54",x"4f"),
  2496 => (x"45",x"4e",x"00",x"53"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

