library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7c40407c",
     1 => x"1c00007c",
     2 => x"3c60603c",
     3 => x"7c3c001c",
     4 => x"7c603060",
     5 => x"6c44003c",
     6 => x"6c381038",
     7 => x"1c000044",
     8 => x"3c60e0bc",
     9 => x"4400001c",
    10 => x"4c5c7464",
    11 => x"08000044",
    12 => x"41773e08",
    13 => x"00000041",
    14 => x"007f7f00",
    15 => x"41000000",
    16 => x"083e7741",
    17 => x"01020008",
    18 => x"02020301",
    19 => x"7f7f0001",
    20 => x"7f7f7f7f",
    21 => x"0808007f",
    22 => x"3e3e1c1c",
    23 => x"7f7f7f7f",
    24 => x"1c1c3e3e",
    25 => x"10000808",
    26 => x"187c7c18",
    27 => x"10000010",
    28 => x"307c7c30",
    29 => x"30100010",
    30 => x"1e786060",
    31 => x"66420006",
    32 => x"663c183c",
    33 => x"38780042",
    34 => x"6cc6c26a",
    35 => x"00600038",
    36 => x"00006000",
    37 => x"5e0e0060",
    38 => x"0e5d5c5b",
    39 => x"c24c711e",
    40 => x"4dbfc5ee",
    41 => x"1ec04bc0",
    42 => x"c702ab74",
    43 => x"48a6c487",
    44 => x"87c578c0",
    45 => x"c148a6c4",
    46 => x"1e66c478",
    47 => x"dfee4973",
    48 => x"c086c887",
    49 => x"efef49e0",
    50 => x"4aa5c487",
    51 => x"f0f0496a",
    52 => x"87c6f187",
    53 => x"83c185cb",
    54 => x"04abb7c8",
    55 => x"2687c7ff",
    56 => x"4c264d26",
    57 => x"4f264b26",
    58 => x"c24a711e",
    59 => x"c25ac9ee",
    60 => x"c748c9ee",
    61 => x"ddfe4978",
    62 => x"1e4f2687",
    63 => x"4a711e73",
    64 => x"03aab7c0",
    65 => x"d2c287d3",
    66 => x"c405bfee",
    67 => x"c24bc187",
    68 => x"c24bc087",
    69 => x"c45bf2d2",
    70 => x"f2d2c287",
    71 => x"eed2c25a",
    72 => x"9ac14abf",
    73 => x"49a2c0c1",
    74 => x"fc87e8ec",
    75 => x"eed2c248",
    76 => x"effe78bf",
    77 => x"4a711e87",
    78 => x"721e66c4",
    79 => x"87f9ea49",
    80 => x"1e4f2626",
    81 => x"d4ff4a71",
    82 => x"78ffc348",
    83 => x"c048d0ff",
    84 => x"d4ff78e1",
    85 => x"7278c148",
    86 => x"7131c449",
    87 => x"48d0ff78",
    88 => x"2678e0c0",
    89 => x"d2c21e4f",
    90 => x"e649bfee",
    91 => x"edc287f9",
    92 => x"bfe848fd",
    93 => x"f9edc278",
    94 => x"78bfec48",
    95 => x"bffdedc2",
    96 => x"ffc3494a",
    97 => x"2ab7c899",
    98 => x"b0714872",
    99 => x"58c5eec2",
   100 => x"5e0e4f26",
   101 => x"0e5d5c5b",
   102 => x"c8ff4b71",
   103 => x"f8edc287",
   104 => x"7350c048",
   105 => x"87dfe649",
   106 => x"c24c4970",
   107 => x"49eecb9c",
   108 => x"7087c3cc",
   109 => x"edc24d49",
   110 => x"05bf97f8",
   111 => x"d087e2c1",
   112 => x"eec24966",
   113 => x"0599bfc1",
   114 => x"66d487d6",
   115 => x"f9edc249",
   116 => x"cb0599bf",
   117 => x"e5497387",
   118 => x"987087ed",
   119 => x"87c1c102",
   120 => x"c0fe4cc1",
   121 => x"cb497587",
   122 => x"987087d8",
   123 => x"c287c602",
   124 => x"c148f8ed",
   125 => x"f8edc250",
   126 => x"c005bf97",
   127 => x"eec287e3",
   128 => x"d049bfc1",
   129 => x"ff059966",
   130 => x"edc287d6",
   131 => x"d449bff9",
   132 => x"ff059966",
   133 => x"497387ca",
   134 => x"7087ece4",
   135 => x"fffe0598",
   136 => x"fa487487",
   137 => x"5e0e87fa",
   138 => x"0e5d5c5b",
   139 => x"4dc086f8",
   140 => x"7ebfec4c",
   141 => x"c248a6c4",
   142 => x"78bfc5ee",
   143 => x"1ec01ec1",
   144 => x"cdfd49c7",
   145 => x"7086c887",
   146 => x"87cd0298",
   147 => x"eafa49ff",
   148 => x"49dac187",
   149 => x"c187f0e3",
   150 => x"f8edc24d",
   151 => x"cf02bf97",
   152 => x"e6d2c287",
   153 => x"b9c149bf",
   154 => x"59ead2c2",
   155 => x"87d3fb71",
   156 => x"bffdedc2",
   157 => x"eed2c24b",
   158 => x"d9c105bf",
   159 => x"48a6c487",
   160 => x"78c0c0c8",
   161 => x"7ee1dbc2",
   162 => x"49bf976e",
   163 => x"80c1486e",
   164 => x"e2717e70",
   165 => x"987087f1",
   166 => x"c487c302",
   167 => x"66c4b366",
   168 => x"28b7c148",
   169 => x"7058a6c8",
   170 => x"dbff0598",
   171 => x"49fdc387",
   172 => x"c387d4e2",
   173 => x"cee249fa",
   174 => x"c3497387",
   175 => x"1e7199ff",
   176 => x"f0f949c0",
   177 => x"c8497387",
   178 => x"1e7129b7",
   179 => x"e4f949c1",
   180 => x"c586c887",
   181 => x"eec287fa",
   182 => x"9b4bbfc1",
   183 => x"c287dd02",
   184 => x"49bfead2",
   185 => x"7087dbc7",
   186 => x"87c40598",
   187 => x"87d24bc0",
   188 => x"c749e0c2",
   189 => x"d2c287c0",
   190 => x"87c658ee",
   191 => x"48ead2c2",
   192 => x"497378c0",
   193 => x"ce0599c2",
   194 => x"49ebc387",
   195 => x"7087f8e0",
   196 => x"0299c249",
   197 => x"fb87c2c0",
   198 => x"c149734c",
   199 => x"87ce0599",
   200 => x"e049f4c3",
   201 => x"497087e1",
   202 => x"c00299c2",
   203 => x"4cfa87c2",
   204 => x"99c84973",
   205 => x"c387cd05",
   206 => x"cae049f5",
   207 => x"c2497087",
   208 => x"87d60299",
   209 => x"bfc9eec2",
   210 => x"87cac002",
   211 => x"c288c148",
   212 => x"c058cdee",
   213 => x"4cff87c2",
   214 => x"49734dc1",
   215 => x"c00599c4",
   216 => x"f2c387ce",
   217 => x"dedfff49",
   218 => x"c2497087",
   219 => x"87dc0299",
   220 => x"bfc9eec2",
   221 => x"b7c7487e",
   222 => x"cbc003a8",
   223 => x"c1486e87",
   224 => x"cdeec280",
   225 => x"87c2c058",
   226 => x"4dc14cfe",
   227 => x"ff49fdc3",
   228 => x"7087f4de",
   229 => x"0299c249",
   230 => x"c287d5c0",
   231 => x"02bfc9ee",
   232 => x"c287c9c0",
   233 => x"c048c9ee",
   234 => x"87c2c078",
   235 => x"4dc14cfd",
   236 => x"ff49fac3",
   237 => x"7087d0de",
   238 => x"0299c249",
   239 => x"c287d9c0",
   240 => x"48bfc9ee",
   241 => x"03a8b7c7",
   242 => x"c287c9c0",
   243 => x"c748c9ee",
   244 => x"87c2c078",
   245 => x"4dc14cfc",
   246 => x"03acb7c0",
   247 => x"c487d3c0",
   248 => x"d8c14866",
   249 => x"6e7e7080",
   250 => x"c5c002bf",
   251 => x"49744b87",
   252 => x"1ec00f73",
   253 => x"c11ef0c3",
   254 => x"d5f649da",
   255 => x"7086c887",
   256 => x"d8c00298",
   257 => x"c9eec287",
   258 => x"496e7ebf",
   259 => x"66c491cb",
   260 => x"6a82714a",
   261 => x"87c5c002",
   262 => x"73496e4b",
   263 => x"029d750f",
   264 => x"c287c8c0",
   265 => x"49bfc9ee",
   266 => x"c287ebf1",
   267 => x"02bff2d2",
   268 => x"4987ddc0",
   269 => x"7087cbc2",
   270 => x"d3c00298",
   271 => x"c9eec287",
   272 => x"d1f149bf",
   273 => x"f249c087",
   274 => x"d2c287f1",
   275 => x"78c048f2",
   276 => x"cbf28ef8",
   277 => x"5b5e0e87",
   278 => x"1e0e5d5c",
   279 => x"eec24c71",
   280 => x"c149bfc5",
   281 => x"c14da1cd",
   282 => x"7e6981d1",
   283 => x"cf029c74",
   284 => x"4ba5c487",
   285 => x"eec27b74",
   286 => x"f149bfc5",
   287 => x"7b6e87ea",
   288 => x"c4059c74",
   289 => x"c24bc087",
   290 => x"734bc187",
   291 => x"87ebf149",
   292 => x"c70266d4",
   293 => x"87de4987",
   294 => x"87c24a70",
   295 => x"d2c24ac0",
   296 => x"f0265af6",
   297 => x"000087fa",
   298 => x"00000000",
   299 => x"00000000",
   300 => x"00000000",
   301 => x"711e0000",
   302 => x"bfc8ff4a",
   303 => x"48a17249",
   304 => x"ff1e4f26",
   305 => x"fe89bfc8",
   306 => x"c0c0c0c0",
   307 => x"c401a9c0",
   308 => x"c24ac087",
   309 => x"724ac187",
   310 => x"0e4f2648",
   311 => x"5d5c5b5e",
   312 => x"ff4b710e",
   313 => x"66d04cd4",
   314 => x"d678c048",
   315 => x"cedbff49",
   316 => x"7cffc387",
   317 => x"ffc3496c",
   318 => x"494d7199",
   319 => x"c199f0c3",
   320 => x"cb05a9e0",
   321 => x"7cffc387",
   322 => x"98c3486c",
   323 => x"780866d0",
   324 => x"6c7cffc3",
   325 => x"31c8494a",
   326 => x"6c7cffc3",
   327 => x"72b2714a",
   328 => x"c331c849",
   329 => x"4a6c7cff",
   330 => x"4972b271",
   331 => x"ffc331c8",
   332 => x"714a6c7c",
   333 => x"48d0ffb2",
   334 => x"7378e0c0",
   335 => x"87c2029b",
   336 => x"48757b72",
   337 => x"4c264d26",
   338 => x"4f264b26",
   339 => x"0e4f261e",
   340 => x"0e5c5b5e",
   341 => x"1e7686f8",
   342 => x"fd49a6c8",
   343 => x"86c487fd",
   344 => x"486e4b70",
   345 => x"c203a8c2",
   346 => x"4a7387f0",
   347 => x"c19af0c3",
   348 => x"c702aad0",
   349 => x"aae0c187",
   350 => x"87dec205",
   351 => x"99c84973",
   352 => x"ff87c302",
   353 => x"4c7387c6",
   354 => x"acc29cc3",
   355 => x"87c2c105",
   356 => x"c94966c4",
   357 => x"c41e7131",
   358 => x"92d44a66",
   359 => x"49cdeec2",
   360 => x"d0fe8172",
   361 => x"49d887eb",
   362 => x"87d3d8ff",
   363 => x"c21ec0c8",
   364 => x"fd49eadc",
   365 => x"ff87e7ec",
   366 => x"e0c048d0",
   367 => x"eadcc278",
   368 => x"4a66cc1e",
   369 => x"eec292d4",
   370 => x"817249cd",
   371 => x"87f2cefe",
   372 => x"acc186cc",
   373 => x"87c2c105",
   374 => x"c94966c4",
   375 => x"c41e7131",
   376 => x"92d44a66",
   377 => x"49cdeec2",
   378 => x"cffe8172",
   379 => x"dcc287e3",
   380 => x"66c81eea",
   381 => x"c292d44a",
   382 => x"7249cdee",
   383 => x"f2ccfe81",
   384 => x"ff49d787",
   385 => x"c887f8d6",
   386 => x"dcc21ec0",
   387 => x"eafd49ea",
   388 => x"86cc87e5",
   389 => x"c048d0ff",
   390 => x"8ef878e0",
   391 => x"0e87e7fc",
   392 => x"5d5c5b5e",
   393 => x"4d711e0e",
   394 => x"d44cd4ff",
   395 => x"c3487e66",
   396 => x"c506a8b7",
   397 => x"c148c087",
   398 => x"497587e2",
   399 => x"87deddfe",
   400 => x"66c41e75",
   401 => x"c293d44b",
   402 => x"7383cdee",
   403 => x"efc6fe49",
   404 => x"6b83c887",
   405 => x"48d0ff4b",
   406 => x"dd78e1c8",
   407 => x"c349737c",
   408 => x"7c7199ff",
   409 => x"b7c84973",
   410 => x"99ffc329",
   411 => x"49737c71",
   412 => x"c329b7d0",
   413 => x"7c7199ff",
   414 => x"b7d84973",
   415 => x"c07c7129",
   416 => x"7c7c7c7c",
   417 => x"7c7c7c7c",
   418 => x"7c7c7c7c",
   419 => x"c478e0c0",
   420 => x"49dc1e66",
   421 => x"87ccd5ff",
   422 => x"487386c8",
   423 => x"87e4fa26",
   424 => x"c01e731e",
   425 => x"f5dbc24b",
   426 => x"c250c048",
   427 => x"49bff1db",
   428 => x"87cedffe",
   429 => x"c4059870",
   430 => x"c9dbc287",
   431 => x"c448734b",
   432 => x"264d2687",
   433 => x"264b264c",
   434 => x"6f68534f",
   435 => x"69682f77",
   436 => x"4f206564",
   437 => x"3d204453",
   438 => x"79656b20",
   439 => x"32314620",
   440 => x"14125800",
   441 => x"1c1b1d11",
   442 => x"94595a23",
   443 => x"ebf2f591",
   444 => x"0026f6f4",
   445 => x"55410000",
   446 => x"4f424f54",
   447 => x"454e544f",
   448 => x"454e0053",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
